-- Version: v11.7 11.7.0.119

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity M2sExt_sb_MSS is

    port( USB_ULPI_DATA                               : inout std_logic_vector(7 downto 0) := (others => 'Z');
          GPOUT_reg                                   : in    std_logic_vector(3 to 3);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR  : inout std_logic_vector(15 downto 12) := (others => 'Z');
          CoreAPB3_0_APBmslave0_PADDR                 : inout std_logic_vector(8 downto 0) := (others => 'Z');
          CoreAPB3_0_APBmslave0_PWDATA                : out   std_logic_vector(31 downto 0);
          COREI2C_0_0_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_1_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_2_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_3_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_4_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_5_INT                             : in    std_logic_vector(0 to 0);
          COREI2C_0_6_INT                             : in    std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : in    std_logic_vector(31 downto 8);
          USB_ULPI_XCLK                               : in    std_logic;
          USB_ULPI_STP                                : out   std_logic;
          USB_ULPI_NXT                                : in    std_logic;
          USB_ULPI_DIR                                : in    std_logic;
          N_48                                        : in    std_logic;
          un561_psel_4                                : in    std_logic;
          m7_x                                        : in    std_logic;
          N_47                                        : in    std_logic;
          N_1217                                      : in    std_logic;
          N_1217_0                                    : in    std_logic;
          N_1217_1                                    : in    std_logic;
          N_1217_2                                    : in    std_logic;
          N_8_0                                       : in    std_logic;
          m71_1                                       : in    std_logic;
          N_1217_3                                    : in    std_logic;
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : inout std_logic := 'Z';
          CoreAPB3_0_APBmslave7_PSELx                 : in    std_logic;
          un30_psel                                   : in    std_logic;
          N_6186                                      : in    std_logic;
          M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N    : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE               : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                : out   std_logic;
          M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F         : out   std_logic;
          N_23_0_i_0                                  : in    std_logic;
          N_38_i_0                                    : in    std_logic;
          N_62_i_0                                    : in    std_logic;
          N_92_i_0                                    : in    std_logic;
          N_107_i_0                                   : in    std_logic;
          N_122_i_0                                   : in    std_logic;
          N_137_i_0                                   : in    std_logic;
          FAB_CCC_LOCK                                : in    std_logic;
          FAB_CCC_GL0                                 : in    std_logic
        );

end M2sExt_sb_MSS;

architecture DEF_ARCH of M2sExt_sb_MSS is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component MSS_010

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic
        );
  end component;

    signal USB_ULPI_XCLK_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE, 
        USB_ULPI_NXT_PAD_Y, USB_ULPI_DIR_PAD_Y, 
        USB_ULPI_DATA_7_PAD_Y, 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, 
        USB_ULPI_DATA_6_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT, 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE, 
        USB_ULPI_DATA_5_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT, 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE, 
        USB_ULPI_DATA_4_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT, 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE, 
        USB_ULPI_DATA_3_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, 
        USB_ULPI_DATA_2_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        USB_ULPI_DATA_1_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, 
        USB_ULPI_DATA_0_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, 
        d_m7_1_0_1, N_6, N_16, G_17_0_1, N_77_i_0, G_17_0_a6_1_4, 
        G_17_0_a6_1_3, G_17_0_1_0, G_17_0_a6_0_1, G_17_0_m6_1, 
        N_9, G_17_0_a6_0_1_1, G_17_0_a6_3_3, VCC_net_1, GND_net_1
         : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc329, 
        nc66, nc83, nc9, nc252, nc171, nc54, nc286, nc307, nc135, 
        nc41, nc100, nc270, nc52, nc251, nc186, nc29, nc269, 
        nc118, nc60, nc141, nc311, nc276, nc193, nc214, nc298, 
        nc282, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc281, nc209, nc246, nc162, nc11, nc272, nc131, nc254, 
        nc267, nc96, nc79, nc226, nc146, nc230, nc89, nc119, nc48, 
        nc271, nc213, nc300, nc126, nc195, nc188, nc242, nc15, 
        nc308, nc236, nc102, nc304, nc3, nc207, nc47, nc90, nc284, 
        nc222, nc159, nc136, nc241, nc253, nc178, nc306, nc215, 
        nc59, nc221, nc232, nc274, nc18, nc44, nc117, nc189, 
        nc164, nc148, nc42, nc231, nc191, nc255, nc283, nc317, 
        nc290, nc17, nc2, nc302, nc110, nc128, nc244, nc321, nc43, 
        nc179, nc157, nc36, nc224, nc296, nc273, nc61, nc104, 
        nc138, nc14, nc285, nc303, nc150, nc196, nc234, nc149, 
        nc12, nc219, nc30, nc243, nc187, nc65, nc7, nc292, nc129, 
        nc275, nc8, nc223, nc13, nc305, nc180, nc26, nc291, nc177, 
        nc139, nc310, nc259, nc245, nc233, nc163, nc318, nc268, 
        nc112, nc68, nc49, nc314, nc217, nc170, nc91, nc225, nc5, 
        nc20, nc198, nc147, nc316, nc67, nc289, nc294, nc152, 
        nc127, nc103, nc235, nc76, nc208, nc140, nc257, nc86, 
        nc95, nc327, nc120, nc165, nc279, nc137, nc64, nc19, 
        nc312, nc70, nc182, nc62, nc199, nc80, nc130, nc287, nc98, 
        nc293, nc249, nc114, nc56, nc105, nc63, nc313, nc309, 
        nc172, nc229, nc277, nc97, nc161, nc31, nc295, nc154, 
        nc50, nc260, nc239, nc142, nc320, nc315, nc247, nc94, 
        nc197, nc328, nc122, nc266, nc35, nc324, nc4, nc227, nc92, 
        nc101, nc330, nc184, nc200, nc190, nc166, nc326, nc132, 
        nc21, nc237, nc93, nc262, nc69, nc206, nc174, nc38, nc113, 
        nc218, nc106, nc261, nc25, nc1, nc322, nc299, nc37, nc202, 
        nc144, nc153, nc46, nc258, nc71, nc124, nc81, nc201, 
        nc168, nc323, nc34, nc28, nc115, nc264, nc192, nc319, 
        nc134, nc32, nc40, nc297, nc99, nc75, nc183, nc288, nc85, 
        nc27, nc108, nc325, nc16, nc155, nc51, nc301, nc33, nc204, 
        nc173, nc278, nc169, nc78, nc263, nc24, nc88, nc111, nc55, 
        nc10, nc22, nc210, nc185, nc143, nc248, nc77, nc6, nc109, 
        nc87, nc123 : std_logic;

begin 


    MSS_ADLIB_INST_RNO_7 : CFG4
      generic map(INIT => x"0040")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        G_17_0_a6_0_1_1, C => N_8_0, D => m71_1, Y => 
        G_17_0_a6_0_1);
    
    MSS_ADLIB_INST_RNO_0 : CFG4
      generic map(INIT => x"FDF5")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => un30_psel, D => 
        N_6186, Y => N_6);
    
    USB_ULPI_DATA_5_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(5), D => 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT, E => 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE, Y => 
        USB_ULPI_DATA_5_PAD_Y);
    
    USB_ULPI_DIR_PAD : INBUF
      port map(PAD => USB_ULPI_DIR, Y => USB_ULPI_DIR_PAD_Y);
    
    USB_ULPI_DATA_2_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(2), D => 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, E
         => MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        Y => USB_ULPI_DATA_2_PAD_Y);
    
    USB_ULPI_DATA_0_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(0), D => 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, E => 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, Y => 
        USB_ULPI_DATA_0_PAD_Y);
    
    MSS_ADLIB_INST_RNO : CFG4
      generic map(INIT => x"DCFE")

      port map(A => N_6, B => N_16, C => N_47, D => G_17_0_1, Y
         => N_77_i_0);
    
    MSS_ADLIB_INST_RNO_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), C => 
        GPOUT_reg(3), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, Y => 
        G_17_0_a6_3_3);
    
    MSS_ADLIB_INST_RNO_5 : CFG3
      generic map(INIT => x"10")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => N_1217_3, Y => 
        G_17_0_a6_1_3);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNO_8 : CFG4
      generic map(INIT => x"A0DD")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1217, C => N_1217_0, D => G_17_0_m6_1, Y => N_9);
    
    USB_ULPI_NXT_PAD : INBUF
      port map(PAD => USB_ULPI_NXT, Y => USB_ULPI_NXT_PAD_Y);
    
    USB_ULPI_DATA_1_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(1), D => 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, E => 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, Y => 
        USB_ULPI_DATA_1_PAD_Y);
    
    USB_ULPI_XCLK_PAD : INBUF
      port map(PAD => USB_ULPI_XCLK, Y => USB_ULPI_XCLK_PAD_Y);
    
    USB_ULPI_DATA_4_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(4), D => 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT, E => 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE, Y => 
        USB_ULPI_DATA_4_PAD_Y);
    
    USB_ULPI_DATA_7_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(7), D => 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, E => 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, Y => 
        USB_ULPI_DATA_7_PAD_Y);
    
    USB_ULPI_STP_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, E => 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE, PAD => 
        USB_ULPI_STP);
    
    MSS_ADLIB_INST_RNO_11 : CFG4
      generic map(INIT => x"2367")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        N_1217_1, D => N_1217_2, Y => G_17_0_m6_1);
    
    USB_ULPI_DATA_3_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(3), D => 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, E
         => MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, Y
         => USB_ULPI_DATA_3_PAD_Y);
    
    MSS_ADLIB_INST_RNO_4 : CFG4
      generic map(INIT => x"8000")

      port map(A => un561_psel_4, B => N_8_0, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), Y => 
        G_17_0_a6_1_4);
    
    MSS_ADLIB_INST_RNO_2 : CFG4
      generic map(INIT => x"0007")

      port map(A => G_17_0_a6_1_4, B => G_17_0_a6_1_3, C => 
        G_17_0_1_0, D => G_17_0_a6_0_1, Y => G_17_0_1);
    
    MSS_ADLIB_INST_RNO_10 : CFG3
      generic map(INIT => x"20")

      port map(A => un561_psel_4, B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), Y => 
        G_17_0_a6_0_1_1);
    
    MSS_ADLIB_INST_RNO_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15), C => 
        un30_psel, D => G_17_0_a6_3_3, Y => N_16);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    USB_ULPI_DATA_6_PAD : BIBUF
      port map(PAD => USB_ULPI_DATA(6), D => 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT, E => 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE, Y => 
        USB_ULPI_DATA_6_PAD_Y);
    
    MSS_ADLIB_INST_RNO_6 : CFG3
      generic map(INIT => x"20")

      port map(A => N_9, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => 
        d_m7_1_0_1, Y => G_17_0_1_0);
    
    MSS_ADLIB_INST_RNO_9 : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => N_48, C
         => un561_psel_4, D => m7_x, Y => d_m7_1_0_1);
    
    MSS_ADLIB_INST : MSS_010

              generic map(INIT => "00" & x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000120481204812048120D8120D8120F00000000F000000000000000000000000000000007FFFFFFFB000001007C33D00809000608EC0000003FFFFE400000000002110000000000F01C000001FECFF4010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 0.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, EDAC_ERROR(7)
         => nc228, EDAC_ERROR(6) => nc203, EDAC_ERROR(5) => nc265, 
        EDAC_ERROR(4) => nc216, EDAC_ERROR(3) => nc194, 
        EDAC_ERROR(2) => nc151, EDAC_ERROR(1) => nc23, 
        EDAC_ERROR(0) => nc175, F_FM0_RDATA(31) => nc250, 
        F_FM0_RDATA(30) => nc58, F_FM0_RDATA(29) => nc116, 
        F_FM0_RDATA(28) => nc74, F_FM0_RDATA(27) => nc133, 
        F_FM0_RDATA(26) => nc238, F_FM0_RDATA(25) => nc167, 
        F_FM0_RDATA(24) => nc84, F_FM0_RDATA(23) => nc39, 
        F_FM0_RDATA(22) => nc72, F_FM0_RDATA(21) => nc256, 
        F_FM0_RDATA(20) => nc212, F_FM0_RDATA(19) => nc205, 
        F_FM0_RDATA(18) => nc82, F_FM0_RDATA(17) => nc145, 
        F_FM0_RDATA(16) => nc181, F_FM0_RDATA(15) => nc160, 
        F_FM0_RDATA(14) => nc57, F_FM0_RDATA(13) => nc156, 
        F_FM0_RDATA(12) => nc280, F_FM0_RDATA(11) => nc125, 
        F_FM0_RDATA(10) => nc211, F_FM0_RDATA(9) => nc73, 
        F_FM0_RDATA(8) => nc107, F_FM0_RDATA(7) => nc329, 
        F_FM0_RDATA(6) => nc66, F_FM0_RDATA(5) => nc83, 
        F_FM0_RDATA(4) => nc9, F_FM0_RDATA(3) => nc252, 
        F_FM0_RDATA(2) => nc171, F_FM0_RDATA(1) => nc54, 
        F_FM0_RDATA(0) => nc286, F_FM0_READYOUT => OPEN, 
        F_FM0_RESP => OPEN, F_HM0_ADDR(31) => nc307, 
        F_HM0_ADDR(30) => nc135, F_HM0_ADDR(29) => nc41, 
        F_HM0_ADDR(28) => nc100, F_HM0_ADDR(27) => nc270, 
        F_HM0_ADDR(26) => nc52, F_HM0_ADDR(25) => nc251, 
        F_HM0_ADDR(24) => nc186, F_HM0_ADDR(23) => nc29, 
        F_HM0_ADDR(22) => nc269, F_HM0_ADDR(21) => nc118, 
        F_HM0_ADDR(20) => nc60, F_HM0_ADDR(19) => nc141, 
        F_HM0_ADDR(18) => nc311, F_HM0_ADDR(17) => nc276, 
        F_HM0_ADDR(16) => nc193, F_HM0_ADDR(15) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15), 
        F_HM0_ADDR(14) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), 
        F_HM0_ADDR(13) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), 
        F_HM0_ADDR(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), 
        F_HM0_ADDR(11) => nc214, F_HM0_ADDR(10) => nc298, 
        F_HM0_ADDR(9) => nc282, F_HM0_ADDR(8) => 
        CoreAPB3_0_APBmslave0_PADDR(8), F_HM0_ADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), F_HM0_ADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), F_HM0_ADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), F_HM0_ADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), F_HM0_ADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), F_HM0_ADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), F_HM0_ADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), F_HM0_ADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), F_HM0_ENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, F_HM0_SEL => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, F_HM0_SIZE(1)
         => nc240, F_HM0_SIZE(0) => nc45, F_HM0_TRANS1 => OPEN, 
        F_HM0_WDATA(31) => CoreAPB3_0_APBmslave0_PWDATA(31), 
        F_HM0_WDATA(30) => CoreAPB3_0_APBmslave0_PWDATA(30), 
        F_HM0_WDATA(29) => CoreAPB3_0_APBmslave0_PWDATA(29), 
        F_HM0_WDATA(28) => CoreAPB3_0_APBmslave0_PWDATA(28), 
        F_HM0_WDATA(27) => CoreAPB3_0_APBmslave0_PWDATA(27), 
        F_HM0_WDATA(26) => CoreAPB3_0_APBmslave0_PWDATA(26), 
        F_HM0_WDATA(25) => CoreAPB3_0_APBmslave0_PWDATA(25), 
        F_HM0_WDATA(24) => CoreAPB3_0_APBmslave0_PWDATA(24), 
        F_HM0_WDATA(23) => CoreAPB3_0_APBmslave0_PWDATA(23), 
        F_HM0_WDATA(22) => CoreAPB3_0_APBmslave0_PWDATA(22), 
        F_HM0_WDATA(21) => CoreAPB3_0_APBmslave0_PWDATA(21), 
        F_HM0_WDATA(20) => CoreAPB3_0_APBmslave0_PWDATA(20), 
        F_HM0_WDATA(19) => CoreAPB3_0_APBmslave0_PWDATA(19), 
        F_HM0_WDATA(18) => CoreAPB3_0_APBmslave0_PWDATA(18), 
        F_HM0_WDATA(17) => CoreAPB3_0_APBmslave0_PWDATA(17), 
        F_HM0_WDATA(16) => CoreAPB3_0_APBmslave0_PWDATA(16), 
        F_HM0_WDATA(15) => CoreAPB3_0_APBmslave0_PWDATA(15), 
        F_HM0_WDATA(14) => CoreAPB3_0_APBmslave0_PWDATA(14), 
        F_HM0_WDATA(13) => CoreAPB3_0_APBmslave0_PWDATA(13), 
        F_HM0_WDATA(12) => CoreAPB3_0_APBmslave0_PWDATA(12), 
        F_HM0_WDATA(11) => CoreAPB3_0_APBmslave0_PWDATA(11), 
        F_HM0_WDATA(10) => CoreAPB3_0_APBmslave0_PWDATA(10), 
        F_HM0_WDATA(9) => CoreAPB3_0_APBmslave0_PWDATA(9), 
        F_HM0_WDATA(8) => CoreAPB3_0_APBmslave0_PWDATA(8), 
        F_HM0_WDATA(7) => CoreAPB3_0_APBmslave0_PWDATA(7), 
        F_HM0_WDATA(6) => CoreAPB3_0_APBmslave0_PWDATA(6), 
        F_HM0_WDATA(5) => CoreAPB3_0_APBmslave0_PWDATA(5), 
        F_HM0_WDATA(4) => CoreAPB3_0_APBmslave0_PWDATA(4), 
        F_HM0_WDATA(3) => CoreAPB3_0_APBmslave0_PWDATA(3), 
        F_HM0_WDATA(2) => CoreAPB3_0_APBmslave0_PWDATA(2), 
        F_HM0_WDATA(1) => CoreAPB3_0_APBmslave0_PWDATA(1), 
        F_HM0_WDATA(0) => CoreAPB3_0_APBmslave0_PWDATA(0), 
        F_HM0_WRITE => CoreAPB3_0_APBmslave0_PWRITE, FAB_CHRGVBUS
         => OPEN, FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc53, FAB_OPMODE(0) => nc121, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc176, FAB_VCONTROL(2) => 
        nc220, FAB_VCONTROL(1) => nc158, FAB_VCONTROL(0) => nc281, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc209, 
        FAB_XCVRSEL(0) => nc246, FAB_XDATAOUT(7) => nc162, 
        FAB_XDATAOUT(6) => nc11, FAB_XDATAOUT(5) => nc272, 
        FAB_XDATAOUT(4) => nc131, FAB_XDATAOUT(3) => nc254, 
        FAB_XDATAOUT(2) => nc267, FAB_XDATAOUT(1) => nc96, 
        FAB_XDATAOUT(0) => nc79, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc226, FIC32_0_MASTER(0) => nc146, 
        FIC32_1_MASTER(1) => nc230, FIC32_1_MASTER(0) => nc89, 
        FPGA_RESET_N => M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        GTX_CLK => OPEN, H2F_INTERRUPT(15) => nc119, 
        H2F_INTERRUPT(14) => nc48, H2F_INTERRUPT(13) => nc271, 
        H2F_INTERRUPT(12) => nc213, H2F_INTERRUPT(11) => nc300, 
        H2F_INTERRUPT(10) => nc126, H2F_INTERRUPT(9) => nc195, 
        H2F_INTERRUPT(8) => nc188, H2F_INTERRUPT(7) => nc242, 
        H2F_INTERRUPT(6) => nc15, H2F_INTERRUPT(5) => nc308, 
        H2F_INTERRUPT(4) => nc236, H2F_INTERRUPT(3) => nc102, 
        H2F_INTERRUPT(2) => nc304, H2F_INTERRUPT(1) => nc3, 
        H2F_INTERRUPT(0) => nc207, H2F_NMI => OPEN, H2FCALIB => 
        OPEN, I2C0_SCL_MGPIO31B_H2F_A => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_B => OPEN, I2C0_SDA_MGPIO30B_H2F_A
         => OPEN, I2C0_SDA_MGPIO30B_H2F_B => OPEN, 
        I2C1_SCL_MGPIO1A_H2F_A => OPEN, I2C1_SCL_MGPIO1A_H2F_B
         => OPEN, I2C1_SDA_MGPIO0A_H2F_A => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_B => OPEN, MDCF => OPEN, MDOENF => 
        OPEN, MDOF => OPEN, MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc47, PER2_FABRIC_PADDR(14) => 
        nc90, PER2_FABRIC_PADDR(13) => nc284, 
        PER2_FABRIC_PADDR(12) => nc222, PER2_FABRIC_PADDR(11) => 
        nc159, PER2_FABRIC_PADDR(10) => nc136, 
        PER2_FABRIC_PADDR(9) => nc241, PER2_FABRIC_PADDR(8) => 
        nc253, PER2_FABRIC_PADDR(7) => nc178, 
        PER2_FABRIC_PADDR(6) => nc306, PER2_FABRIC_PADDR(5) => 
        nc215, PER2_FABRIC_PADDR(4) => nc59, PER2_FABRIC_PADDR(3)
         => nc221, PER2_FABRIC_PADDR(2) => nc232, 
        PER2_FABRIC_PENABLE => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc274, PER2_FABRIC_PWDATA(30)
         => nc18, PER2_FABRIC_PWDATA(29) => nc44, 
        PER2_FABRIC_PWDATA(28) => nc117, PER2_FABRIC_PWDATA(27)
         => nc189, PER2_FABRIC_PWDATA(26) => nc164, 
        PER2_FABRIC_PWDATA(25) => nc148, PER2_FABRIC_PWDATA(24)
         => nc42, PER2_FABRIC_PWDATA(23) => nc231, 
        PER2_FABRIC_PWDATA(22) => nc191, PER2_FABRIC_PWDATA(21)
         => nc255, PER2_FABRIC_PWDATA(20) => nc283, 
        PER2_FABRIC_PWDATA(19) => nc317, PER2_FABRIC_PWDATA(18)
         => nc290, PER2_FABRIC_PWDATA(17) => nc17, 
        PER2_FABRIC_PWDATA(16) => nc2, PER2_FABRIC_PWDATA(15) => 
        nc302, PER2_FABRIC_PWDATA(14) => nc110, 
        PER2_FABRIC_PWDATA(13) => nc128, PER2_FABRIC_PWDATA(12)
         => nc244, PER2_FABRIC_PWDATA(11) => nc321, 
        PER2_FABRIC_PWDATA(10) => nc43, PER2_FABRIC_PWDATA(9) => 
        nc179, PER2_FABRIC_PWDATA(8) => nc157, 
        PER2_FABRIC_PWDATA(7) => nc36, PER2_FABRIC_PWDATA(6) => 
        nc224, PER2_FABRIC_PWDATA(5) => nc296, 
        PER2_FABRIC_PWDATA(4) => nc273, PER2_FABRIC_PWDATA(3) => 
        nc61, PER2_FABRIC_PWDATA(2) => nc104, 
        PER2_FABRIC_PWDATA(1) => nc138, PER2_FABRIC_PWDATA(0) => 
        nc14, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => OPEN, SPI1_SDO_MGPIO12A_H2F_A => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_B => OPEN, SPI1_SS0_MGPIO13A_H2F_A
         => OPEN, SPI1_SS0_MGPIO13A_H2F_B => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc285, 
        TCGF(8) => nc303, TCGF(7) => nc150, TCGF(6) => nc196, 
        TCGF(5) => nc234, TCGF(4) => nc149, TCGF(3) => nc12, 
        TCGF(2) => nc219, TCGF(1) => nc30, TCGF(0) => nc243, 
        TRACECLK => OPEN, TRACEDATA(3) => nc187, TRACEDATA(2) => 
        nc65, TRACEDATA(1) => nc7, TRACEDATA(0) => nc292, TX_CLK
         => OPEN, TX_ENF => OPEN, TX_ERRF => OPEN, TXCTL_EN_RIF
         => OPEN, TXD_RIF(3) => nc129, TXD_RIF(2) => nc275, 
        TXD_RIF(1) => nc8, TXD_RIF(0) => nc223, TXDF(7) => nc13, 
        TXDF(6) => nc305, TXDF(5) => nc180, TXDF(4) => nc26, 
        TXDF(3) => nc291, TXDF(2) => nc177, TXDF(1) => nc139, 
        TXDF(0) => nc310, TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc259, F_BID(2) => nc245, F_BID(1) => 
        nc233, F_BID(0) => nc163, F_BRESP_HRESP0(1) => nc318, 
        F_BRESP_HRESP0(0) => nc268, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc112, F_RDATA_HRDATA01(62) => 
        nc68, F_RDATA_HRDATA01(61) => nc49, F_RDATA_HRDATA01(60)
         => nc314, F_RDATA_HRDATA01(59) => nc217, 
        F_RDATA_HRDATA01(58) => nc170, F_RDATA_HRDATA01(57) => 
        nc91, F_RDATA_HRDATA01(56) => nc225, F_RDATA_HRDATA01(55)
         => nc5, F_RDATA_HRDATA01(54) => nc20, 
        F_RDATA_HRDATA01(53) => nc198, F_RDATA_HRDATA01(52) => 
        nc147, F_RDATA_HRDATA01(51) => nc316, 
        F_RDATA_HRDATA01(50) => nc67, F_RDATA_HRDATA01(49) => 
        nc289, F_RDATA_HRDATA01(48) => nc294, 
        F_RDATA_HRDATA01(47) => nc152, F_RDATA_HRDATA01(46) => 
        nc127, F_RDATA_HRDATA01(45) => nc103, 
        F_RDATA_HRDATA01(44) => nc235, F_RDATA_HRDATA01(43) => 
        nc76, F_RDATA_HRDATA01(42) => nc208, F_RDATA_HRDATA01(41)
         => nc140, F_RDATA_HRDATA01(40) => nc257, 
        F_RDATA_HRDATA01(39) => nc86, F_RDATA_HRDATA01(38) => 
        nc95, F_RDATA_HRDATA01(37) => nc327, F_RDATA_HRDATA01(36)
         => nc120, F_RDATA_HRDATA01(35) => nc165, 
        F_RDATA_HRDATA01(34) => nc279, F_RDATA_HRDATA01(33) => 
        nc137, F_RDATA_HRDATA01(32) => nc64, F_RDATA_HRDATA01(31)
         => nc19, F_RDATA_HRDATA01(30) => nc312, 
        F_RDATA_HRDATA01(29) => nc70, F_RDATA_HRDATA01(28) => 
        nc182, F_RDATA_HRDATA01(27) => nc62, F_RDATA_HRDATA01(26)
         => nc199, F_RDATA_HRDATA01(25) => nc80, 
        F_RDATA_HRDATA01(24) => nc130, F_RDATA_HRDATA01(23) => 
        nc287, F_RDATA_HRDATA01(22) => nc98, F_RDATA_HRDATA01(21)
         => nc293, F_RDATA_HRDATA01(20) => nc249, 
        F_RDATA_HRDATA01(19) => nc114, F_RDATA_HRDATA01(18) => 
        nc56, F_RDATA_HRDATA01(17) => nc105, F_RDATA_HRDATA01(16)
         => nc63, F_RDATA_HRDATA01(15) => nc313, 
        F_RDATA_HRDATA01(14) => nc309, F_RDATA_HRDATA01(13) => 
        nc172, F_RDATA_HRDATA01(12) => nc229, 
        F_RDATA_HRDATA01(11) => nc277, F_RDATA_HRDATA01(10) => 
        nc97, F_RDATA_HRDATA01(9) => nc161, F_RDATA_HRDATA01(8)
         => nc31, F_RDATA_HRDATA01(7) => nc295, 
        F_RDATA_HRDATA01(6) => nc154, F_RDATA_HRDATA01(5) => nc50, 
        F_RDATA_HRDATA01(4) => nc260, F_RDATA_HRDATA01(3) => 
        nc239, F_RDATA_HRDATA01(2) => nc142, F_RDATA_HRDATA01(1)
         => nc320, F_RDATA_HRDATA01(0) => nc315, F_RID(3) => 
        nc247, F_RID(2) => nc94, F_RID(1) => nc197, F_RID(0) => 
        nc328, F_RLAST => OPEN, F_RRESP_HRESP1(1) => nc122, 
        F_RRESP_HRESP1(0) => nc266, F_RVALID => OPEN, F_WREADY
         => OPEN, MDDR_FABRIC_PRDATA(15) => nc35, 
        MDDR_FABRIC_PRDATA(14) => nc324, MDDR_FABRIC_PRDATA(13)
         => nc4, MDDR_FABRIC_PRDATA(12) => nc227, 
        MDDR_FABRIC_PRDATA(11) => nc92, MDDR_FABRIC_PRDATA(10)
         => nc101, MDDR_FABRIC_PRDATA(9) => nc330, 
        MDDR_FABRIC_PRDATA(8) => nc184, MDDR_FABRIC_PRDATA(7) => 
        nc200, MDDR_FABRIC_PRDATA(6) => nc190, 
        MDDR_FABRIC_PRDATA(5) => nc166, MDDR_FABRIC_PRDATA(4) => 
        nc326, MDDR_FABRIC_PRDATA(3) => nc132, 
        MDDR_FABRIC_PRDATA(2) => nc21, MDDR_FABRIC_PRDATA(1) => 
        nc237, MDDR_FABRIC_PRDATA(0) => nc93, MDDR_FABRIC_PREADY
         => OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        COREI2C_0_6_INT(0), F2H_INTERRUPT(5) => 
        COREI2C_0_5_INT(0), F2H_INTERRUPT(4) => 
        COREI2C_0_4_INT(0), F2H_INTERRUPT(3) => 
        COREI2C_0_3_INT(0), F2H_INTERRUPT(2) => 
        COREI2C_0_2_INT(0), F2H_INTERRUPT(1) => 
        COREI2C_0_1_INT(0), F2H_INTERRUPT(0) => 
        COREI2C_0_0_INT(0), F2HCALIB => VCC_net_1, F_DMAREADY(1)
         => VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31)
         => GND_net_1, F_FM0_ADDR(30) => GND_net_1, 
        F_FM0_ADDR(29) => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        F_HM0_RDATA(30) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        F_HM0_RDATA(29) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        F_HM0_RDATA(28) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        F_HM0_RDATA(27) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        F_HM0_RDATA(26) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        F_HM0_RDATA(25) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        F_HM0_RDATA(24) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        F_HM0_RDATA(23) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        F_HM0_RDATA(22) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        F_HM0_RDATA(21) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        F_HM0_RDATA(20) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        F_HM0_RDATA(19) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        F_HM0_RDATA(18) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        F_HM0_RDATA(17) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        F_HM0_RDATA(16) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        F_HM0_RDATA(15) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        F_HM0_RDATA(14) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        F_HM0_RDATA(13) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        F_HM0_RDATA(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        F_HM0_RDATA(11) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        F_HM0_RDATA(10) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        F_HM0_RDATA(9) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        F_HM0_RDATA(8) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        F_HM0_RDATA(7) => N_137_i_0, F_HM0_RDATA(6) => N_122_i_0, 
        F_HM0_RDATA(5) => N_107_i_0, F_HM0_RDATA(4) => N_92_i_0, 
        F_HM0_RDATA(3) => N_77_i_0, F_HM0_RDATA(2) => N_62_i_0, 
        F_HM0_RDATA(1) => N_38_i_0, F_HM0_RDATA(0) => N_23_0_i_0, 
        F_HM0_READY => VCC_net_1, F_HM0_RESP => GND_net_1, 
        FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => VCC_net_1, 
        FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => VCC_net_1, 
        FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N => 
        VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE => 
        VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => VCC_net_1, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => VCC_net_1, 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => VCC_net_1, MGPIO1A_F2H_GPIN => 
        VCC_net_1, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => VCC_net_1, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        VCC_net_1, MGPIO2A_F2H_GPIN => VCC_net_1, 
        MGPIO30B_F2H_GPIN => VCC_net_1, MGPIO31B_F2H_GPIN => 
        VCC_net_1, MGPIO3A_F2H_GPIN => VCC_net_1, 
        MGPIO4A_F2H_GPIN => VCC_net_1, MGPIO5A_F2H_GPIN => 
        VCC_net_1, MGPIO6A_F2H_GPIN => VCC_net_1, 
        MGPIO7A_F2H_GPIN => VCC_net_1, MGPIO8A_F2H_GPIN => 
        VCC_net_1, MGPIO9A_F2H_GPIN => VCC_net_1, 
        MMUART0_CTS_F2H_SCP => VCC_net_1, MMUART0_DCD_F2H_SCP => 
        VCC_net_1, MMUART0_DSR_F2H_SCP => VCC_net_1, 
        MMUART0_DTR_F2H_SCP => VCC_net_1, MMUART0_RI_F2H_SCP => 
        VCC_net_1, MMUART0_RTS_F2H_SCP => VCC_net_1, 
        MMUART0_RXD_F2H_SCP => VCC_net_1, MMUART0_SCK_F2H_SCP => 
        VCC_net_1, MMUART0_TXD_F2H_SCP => VCC_net_1, 
        MMUART1_CTS_F2H_SCP => VCC_net_1, MMUART1_DCD_F2H_SCP => 
        VCC_net_1, MMUART1_DSR_F2H_SCP => VCC_net_1, 
        MMUART1_RI_F2H_SCP => VCC_net_1, MMUART1_RTS_F2H_SCP => 
        VCC_net_1, MMUART1_RXD_F2H_SCP => VCC_net_1, 
        MMUART1_SCK_F2H_SCP => VCC_net_1, MMUART1_TXD_F2H_SCP => 
        VCC_net_1, PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => FAB_CCC_GL0, CLK_MDDR_APB => VCC_net_1, 
        F_ARADDR_HADDR1(31) => VCC_net_1, F_ARADDR_HADDR1(30) => 
        VCC_net_1, F_ARADDR_HADDR1(29) => VCC_net_1, 
        F_ARADDR_HADDR1(28) => VCC_net_1, F_ARADDR_HADDR1(27) => 
        VCC_net_1, F_ARADDR_HADDR1(26) => VCC_net_1, 
        F_ARADDR_HADDR1(25) => VCC_net_1, F_ARADDR_HADDR1(24) => 
        VCC_net_1, F_ARADDR_HADDR1(23) => VCC_net_1, 
        F_ARADDR_HADDR1(22) => VCC_net_1, F_ARADDR_HADDR1(21) => 
        VCC_net_1, F_ARADDR_HADDR1(20) => VCC_net_1, 
        F_ARADDR_HADDR1(19) => VCC_net_1, F_ARADDR_HADDR1(18) => 
        VCC_net_1, F_ARADDR_HADDR1(17) => VCC_net_1, 
        F_ARADDR_HADDR1(16) => VCC_net_1, F_ARADDR_HADDR1(15) => 
        VCC_net_1, F_ARADDR_HADDR1(14) => VCC_net_1, 
        F_ARADDR_HADDR1(13) => VCC_net_1, F_ARADDR_HADDR1(12) => 
        VCC_net_1, F_ARADDR_HADDR1(11) => VCC_net_1, 
        F_ARADDR_HADDR1(10) => VCC_net_1, F_ARADDR_HADDR1(9) => 
        VCC_net_1, F_ARADDR_HADDR1(8) => VCC_net_1, 
        F_ARADDR_HADDR1(7) => VCC_net_1, F_ARADDR_HADDR1(6) => 
        VCC_net_1, F_ARADDR_HADDR1(5) => VCC_net_1, 
        F_ARADDR_HADDR1(4) => VCC_net_1, F_ARADDR_HADDR1(3) => 
        VCC_net_1, F_ARADDR_HADDR1(2) => VCC_net_1, 
        F_ARADDR_HADDR1(1) => VCC_net_1, F_ARADDR_HADDR1(0) => 
        VCC_net_1, F_ARBURST_HTRANS1(1) => GND_net_1, 
        F_ARBURST_HTRANS1(0) => GND_net_1, F_ARID_HSEL1(3) => 
        GND_net_1, F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1)
         => GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GND_net_1, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => GND_net_1, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => GND_net_1, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => GND_net_1, 
        MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => GND_net_1, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => 
        USB_ULPI_XCLK_PAD_Y, RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => 
        USB_ULPI_DATA_7_PAD_Y, RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => 
        USB_ULPI_DATA_2_PAD_Y, RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN
         => USB_ULPI_DATA_0_PAD_Y, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => 
        USB_ULPI_DATA_1_PAD_Y, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => 
        USB_ULPI_DATA_3_PAD_Y, RGMII_RXD3_USBB_DATA4_IN => 
        USB_ULPI_DATA_4_PAD_Y, RGMII_TX_CLK_IN => GND_net_1, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => USB_ULPI_NXT_PAD_Y, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => USB_ULPI_DIR_PAD_Y, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => USB_ULPI_DATA_5_PAD_Y, 
        RGMII_TXD3_USBB_DATA6_IN => USB_ULPI_DATA_6_PAD_Y, 
        SPI0_SCK_USBA_XCLK_IN => GND_net_1, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => GND_net_1, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => GND_net_1, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, SPI1_SCK_IN
         => GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => GND_net_1, 
        SPI1_SS5_MGPIO18A_IN => GND_net_1, SPI1_SS6_MGPIO23A_IN
         => GND_net_1, SPI1_SS7_MGPIO24A_IN => GND_net_1, 
        USBC_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc262, DRAM_ADDR(14) => nc69, DRAM_ADDR(13) => nc206, 
        DRAM_ADDR(12) => nc174, DRAM_ADDR(11) => nc38, 
        DRAM_ADDR(10) => nc113, DRAM_ADDR(9) => nc218, 
        DRAM_ADDR(8) => nc106, DRAM_ADDR(7) => nc261, 
        DRAM_ADDR(6) => nc25, DRAM_ADDR(5) => nc1, DRAM_ADDR(4)
         => nc322, DRAM_ADDR(3) => nc299, DRAM_ADDR(2) => nc37, 
        DRAM_ADDR(1) => nc202, DRAM_ADDR(0) => nc144, DRAM_BA(2)
         => nc153, DRAM_BA(1) => nc46, DRAM_BA(0) => nc258, 
        DRAM_CASN => OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, 
        DRAM_CSN => OPEN, DRAM_DM_RDQS_OUT(2) => nc71, 
        DRAM_DM_RDQS_OUT(1) => nc124, DRAM_DM_RDQS_OUT(0) => nc81, 
        DRAM_DQ_OUT(17) => nc201, DRAM_DQ_OUT(16) => nc168, 
        DRAM_DQ_OUT(15) => nc323, DRAM_DQ_OUT(14) => nc34, 
        DRAM_DQ_OUT(13) => nc28, DRAM_DQ_OUT(12) => nc115, 
        DRAM_DQ_OUT(11) => nc264, DRAM_DQ_OUT(10) => nc192, 
        DRAM_DQ_OUT(9) => nc319, DRAM_DQ_OUT(8) => nc134, 
        DRAM_DQ_OUT(7) => nc32, DRAM_DQ_OUT(6) => nc40, 
        DRAM_DQ_OUT(5) => nc297, DRAM_DQ_OUT(4) => nc99, 
        DRAM_DQ_OUT(3) => nc75, DRAM_DQ_OUT(2) => nc183, 
        DRAM_DQ_OUT(1) => nc288, DRAM_DQ_OUT(0) => nc85, 
        DRAM_DQS_OUT(2) => nc27, DRAM_DQS_OUT(1) => nc108, 
        DRAM_DQS_OUT(0) => nc325, DRAM_FIFO_WE_OUT(1) => nc16, 
        DRAM_FIFO_WE_OUT(0) => nc155, DRAM_ODT => OPEN, DRAM_RASN
         => OPEN, DRAM_RSTN => OPEN, DRAM_WEN => OPEN, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, 
        RGMII_RXD3_USBB_DATA4_OUT => 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT, 
        RGMII_TX_CLK_OUT => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, 
        RGMII_TXD2_USBB_DATA5_OUT => 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT, 
        RGMII_TXD3_USBB_DATA6_OUT => 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT, 
        SPI0_SCK_USBA_XCLK_OUT => OPEN, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, SPI1_SCK_OUT
         => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => OPEN, 
        SPI1_SS5_MGPIO18A_OUT => OPEN, SPI1_SS6_MGPIO23A_OUT => 
        OPEN, SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => 
        OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc51, 
        DM_OE(1) => nc301, DM_OE(0) => nc33, DRAM_DQ_OE(17) => 
        nc204, DRAM_DQ_OE(16) => nc173, DRAM_DQ_OE(15) => nc278, 
        DRAM_DQ_OE(14) => nc169, DRAM_DQ_OE(13) => nc78, 
        DRAM_DQ_OE(12) => nc263, DRAM_DQ_OE(11) => nc24, 
        DRAM_DQ_OE(10) => nc88, DRAM_DQ_OE(9) => nc111, 
        DRAM_DQ_OE(8) => nc55, DRAM_DQ_OE(7) => nc10, 
        DRAM_DQ_OE(6) => nc22, DRAM_DQ_OE(5) => nc210, 
        DRAM_DQ_OE(4) => nc185, DRAM_DQ_OE(3) => nc143, 
        DRAM_DQ_OE(2) => nc248, DRAM_DQ_OE(1) => nc77, 
        DRAM_DQ_OE(0) => nc6, DRAM_DQS_OE(2) => nc109, 
        DRAM_DQS_OE(1) => nc87, DRAM_DQS_OE(0) => nc123, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, 
        RGMII_RXD3_USBB_DATA4_OE => 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE, RGMII_TX_CLK_OE
         => OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE, 
        RGMII_TXD2_USBB_DATA5_OE => 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE, 
        RGMII_TXD3_USBB_DATA6_OE => 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE, 
        SPI0_SCK_USBA_XCLK_OE => OPEN, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, SPI1_SCK_OE => 
        OPEN, SPI1_SDI_MGPIO11A_OE => OPEN, SPI1_SDO_MGPIO12A_OE
         => OPEN, SPI1_SS0_MGPIO13A_OE => OPEN, 
        SPI1_SS1_MGPIO14A_OE => OPEN, SPI1_SS2_MGPIO15A_OE => 
        OPEN, SPI1_SS3_MGPIO16A_OE => OPEN, SPI1_SS4_MGPIO17A_OE
         => OPEN, SPI1_SS5_MGPIO18A_OE => OPEN, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_2 is

    port( COREI2C_0_3_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          seradr0apb                   : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          N_1217                       : out   std_logic;
          N_1218                       : out   std_logic;
          N_1220                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1221                       : out   std_logic;
          BIBUF_COREI2C_0_3_SDA_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_3_SCL_IO_Y   : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          bclke                        : in    std_logic;
          N_40                         : in    std_logic;
          un3_penable_1                : in    std_logic;
          un105_ens1_1                 : in    std_logic;
          un5_penable_1                : in    std_logic
        );

end COREI2CREAL_6_2;

architecture DEF_ARCH of COREI2CREAL_6_2 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_3_SDAO[0]\, \COREI2C_0_3_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_3_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        un1_serdat_2_sqmuxa_2, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, N_1665, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, N_1470, \ack\, ack_7, N_1449, 
        SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, bsd7_tmp_6, \bsd7\, 
        bsd7_9_iv_i_0, \adrcomp\, N_2176_i_0, 
        adrcomp_2_sqmuxa_i_0_2, \PCLKint\, PCLKint_3, 
        un1_pclkint4_i_0, \ack_bit\, \ack_bit_1_sqmuxa\, 
        \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_2, un1_rtn_3_2, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, PCLK_count2_ov_6_1, 
        \un1_PCLK_count1_0_sqmuxa\, CO1, un13_adrcompen, 
        \adrcomp_2_sqmuxa_i_a2_1_5\, N_2187, N_997, un70_fsmsta, 
        N_1046, \adrcomp_2_sqmuxa_i_o2_1_3\, un16_fsmmod, 
        \sersta_32_5[2]\, N_1586_1, N_2181, N_2177, N_2173_i_1, 
        N_133, un1_fsmmod, N_36_i_1, un136_framesync, N_2196, 
        N_2186, \un1_PCLK_count1_0_sqmuxa_1\, 
        \un1_PCLK_count1_0_sqmuxa_0\, 
        \un1_PCLK_count1_0_sqmuxa_1_0\, CO2, ANC2, N_1002, 
        N_976_i_1, N_68, \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, 
        \fsmsta_cnst[0]\, fsmsta_8_9_509_0_1, N_1717, 
        fsmsta_8_9_509_0, N_1652, fsmsta_8_3_601_0_1, 
        fsmsta_8_3_601_0, \un1_pclk_count1_ov_1_1\, 
        \un1_pclk_count1_ov_1\, \PRDATA_3_1_1[3]\, 
        \PRDATA_3_1_1[4]\, \PRDATA_3_1_1[6]\, \PRDATA_3_1_1[5]\, 
        \PRDATA_3_1_1[7]\, \fsmsta_8_ns_1[29]\, 
        \fsmsta_8_ns_1[28]\, \fsmsta_8_ns_1[16]\, un137_framesync, 
        \fsmsta_8_ns_1[18]\, bsd7_tmp_6_ns_1, bsd7_tmp_6_am_0, 
        un105_ens1, un57_fsmsta, \framesync_7_enl_bm[3]\, 
        \framesync_7_enl_am[3]\, framesync_7_e2, N_2171, 
        \fsmsta_8_0_a2_1[7]\, N_2179, N_161_2, 
        fsmsta_8_5_555_a3_0_2, fsmsta_8_5_555_a3_2, 
        bsd7_tmp_6_sn_m6_0, PCLK_count2_ov_6_0_a2_1_0, 
        \fsmsta_nxt_9_m_0[26]\, \fsmsta_nxt_9_m_0[27]\, 
        un111_fsmdet_0, \sersta_32_i_a2_5[3]\, 
        \adrcomp_2_sqmuxa_i_a3_2\, un139_ens1_0, 
        \adrcomp_2_sqmuxa_i_o2_1_1\, \un1_fsmsta_1_i_0_o2_0\, 
        un135_ens1_2, mst, N_127, N_2178, N_145_2, 
        \un151_framesync\, N_67, N_23, N_64, N_26, 
        un26_adrcompen_3, N_1196, N_1197, N_1198, 
        \serdat_i_m_1[7]\, bsd7_tmp_i_m_1, SDAO_int_7_0_275_1, 
        \adrcomp_2_sqmuxa_i_a3_2_0\, un141_ens1_2, 
        fsmsta_8_28_307_a3_0_0, \SDAO_int_1_sqmuxa_3\, 
        \adrcomp_2_sqmuxa_i_a2_1_2\, \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_10_476_i_a6_1, 
        \fsmmod_ns_i_a4_1_0[2]_net_1\, \sersta_32_4[0]\, 
        \sersta_32_3[0]\, \sersta_32_5[1]\, \sersta_32_4[1]\, 
        fsmsta_8_20_379_i_0_a3_5, fsmsta_8_20_379_i_0_a3_4, 
        \sersta_32_i_a2_7[4]\, \sersta_32_i_a2_6[4]\, 
        \sersta_32_4[2]\, un135_ens1_5, un135_ens1_4, 
        un135_ens1_3, un25_fsmsta_1, \sersta_32_i_a2_8[3]\, 
        \sersta_32_i_a2_7[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, un13_adrcompen_4, 
        m7_5, m7_4, \PCLK_count1_ov_1_sqmuxa_1\, un33_fsmsta, 
        un12_pclk_count1, N_1064, framesync_7_sm0, 
        PCLK_count2_ov_6_0_a2_1_4_tz, N_1040, N_1049, N_1034, 
        N_76, CO1_0, CO2_0, CO1_1, N_117_1, \un1_pclk_count1_ov\, 
        \adrcomp_2_sqmuxa_i_a3_3\, SDAO_int_7_0_275_a5_1, 
        \fsmmod_ns_i_0[2]_net_1\, fsmsta_8_10_476_i_0, 
        \SDAO_int_1_sqmuxa_4\, \adrcomp_2_sqmuxa_i_a2_1_4\, 
        PCLK_count2_ov_6_0_a2_1_3, \adrcomp_2_sqmuxa_i_0_0_0\, 
        \sercon_8_2[4]\, \sersta_32_i_a2_9[4]\, \sersta_32_7[2]\, 
        \sersta_32_i_a2_10[3]\, N_2192, 
        fsmsta_nxt_1_sqmuxa_18_s5_1, un25_fsmsta, 
        fsmsta_nxt_1_sqmuxa_24_s4_1, un19_framesync, 
        un25_framesync, \PCLK_count1_0_sqmuxa_4\, N_104, 
        un74_ens1, N_1656, N_2193, N_191, N_154, un91_ens1, 
        \un1_fsmsta_6\, N_155, N_84, N_63, N_130, N_1041, 
        \un1_pclk_count191\, N_1622_2, N_134, N_120, N_124, N_121, 
        fsmsta_8_3_601_a4_0, fsmsta_8_9_509_a4_0, 
        \SDAO_int_1_sqmuxa_7\, N_1054, \fsmsta_nxt_9_m[22]\, 
        \fsmsta_nxt_9_m[21]\, un115_fsmdet, N_157, N_165, 
        un135_ens1, N_163, \fsmmod_ns_0_a4_0_4[3]_net_1\, N_1060, 
        N_1048, N_126, \PCLK_count1_0_sqmuxa_3\, N_70, N_1624, 
        \fsmsta_8_i_0[25]\, N_80, N_82, fsmsta_8_20_379_i_0_o2_0, 
        \sercon_8_0_1[3]\, \fsmsync_ns_0_0_1[0]_net_1\, 
        fsmsta_8_23_351_i_0_1, \un1_ens1_pre_1_sqmuxa_0_a2_1\, 
        N_1058, N_1465, N_166, N_145, un3_penable, 
        \fsmsync_ns_i_0_1_tz[3]_net_1\, N_1059_1, un92_fsmsta, 
        un1_fsmsta_10_i_0, N_86, N_2199, \PWDATA_i_m_1[7]\, 
        \sercon_8_0_2[3]\, fsmsta_8_2_647_i_0_0, N_1051, N_1486, 
        un134_fsmsta, \serdat_0_sqmuxa\, \framesync_7_m2[3]\, 
        N_161, N_1466, N_152, bsd7_9_iv_1, \serdat_2_sqmuxa\, 
        \un1_serdat40\, \un1_bsd7_1_sqmuxa[0]_net_1\, bsd7_9_iv_2, 
        \serdat_1_sqmuxa_1\, \un1_counter_rst_3\, 
        \un1_serdat_2_sqmuxa_1\ : std_logic;

begin 

    COREI2C_0_3_INT(0) <= \COREI2C_0_3_INT[0]\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \un151_framesync\, B => N_2177, C => N_191, Y
         => un1_fsmsta_10_i_0);
    
    \un1_bsd7_1_sqmuxa[0]\ : CFG4
      generic map(INIT => x"A111")

      port map(A => \COREI2C_0_3_INT[0]\, B => \nedetect\, C => 
        un3_penable, D => un105_ens1_1, Y => 
        \un1_bsd7_1_sqmuxa[0]_net_1\);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    SCLO_int_RNIA863 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_3_SCLO[0]\, Y => 
        COREI2C_0_3_SCLO_i(0));
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_0_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_26, B => \adrcompen\, Y => 
        fsmsta_8_28_307_a3_0_0);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_145_2, 
        Y => N_2171);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_191, B => \un1_fsmsta_6\, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => N_166);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \framesync_7_enl_bm[3]\, B => 
        \framesync_7_enl_am[3]\, C => framesync_7_e2, Y => 
        \framesync_7[3]\);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[2]_net_1\, B => seradr0apb(3), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_3, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_2, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \fsmsync_ns_0_0_a2_2_1[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmmod[4]_net_1\, Y => N_117_1);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_1);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \fsmmod_RNIEQCE1[0]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmmod[5]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        N_1622_2);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns\ : CFG4
      generic map(INIT => x"5404")

      port map(A => \fsmdet[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => bsd7_tmp_6_ns_1, D
         => bsd7_tmp_6_am_0, Y => bsd7_tmp_6);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => un25_fsmsta_1, 
        C => \fsmsta[18]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        un25_fsmsta);
    
    \fsmmod_ns_0_a4_0[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => 
        N_1059_1, Y => N_1051);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sersta_32_5[2]\, B => \sersta_32_7[2]\, C
         => un135_ens1_2, D => \un1_fsmsta_1_i_0_o2_0\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1041, B => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, 
        C => N_1040, Y => \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    un7_fsmsta_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[22]_net_1\, 
        Y => N_2178);
    
    \fsmmod_ns_0[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_1064, B => N_1049, C => un115_fsmdet, D => 
        N_1048, Y => \fsmmod_ns[0]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG3
      generic map(INIT => x"F8")

      port map(A => SDAO_int_7_0_275_a5_1, B => N_1466, C => 
        SDAO_int_7_0_275_1, Y => N_1449);
    
    \sersta_RNIMF942[1]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[4]\, C => \sersta[1]_net_1\, D => 
        seradr0apb(4), Y => N_1218);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_am_RNO\ : CFG2
      generic map(INIT => x"4")

      port map(A => \COREI2C_0_3_INT[0]\, B => \nedetect\, Y => 
        bsd7_tmp_6_sn_m6_0);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \sercon[7]_net_1\, D => 
        \un1_pclk_count1_ov_1_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => un139_ens1_0, Y => 
        framesync_7_sm0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_121, B => N_2181, C => N_154, D => N_155, Y
         => N_2172_i_0);
    
    \fsmmod_ns_0_a4_0[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[1]_net_1\, B => \SCLSCL\, C => 
        \pedetect\, Y => N_1049);
    
    un1_PCLK_count1_0_sqmuxa_0 : CFG4
      generic map(INIT => x"FF10")

      port map(A => \sercon[1]_net_1\, B => \sercon[7]_net_1\, C
         => un12_pclk_count1, D => \PCLK_count1_0_sqmuxa_4\, Y
         => \un1_PCLK_count1_0_sqmuxa_0\);
    
    \fsmsta_RNO[25]\ : CFG3
      generic map(INIT => x"01")

      port map(A => un136_framesync, B => N_154, C => 
        \fsmsta_8_i_0[25]\, Y => N_2175_i_0);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_2_0\, Y
         => \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \fsmsta[17]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_2[3]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \sercon[6]_net_1\, B => \adrcomp\, C => 
        N_1586_1, D => un74_ens1, Y => N_163);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1652, D => un1_fsmmod, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_3_601_0_1);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns_1\ : CFG3
      generic map(INIT => x"7F")

      port map(A => un105_ens1, B => \COREI2C_0_3_INT[0]\, C => 
        un57_fsmsta, Y => bsd7_tmp_6_ns_1);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \serdat_RNIB7DU[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_3_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \serCON_WRITE_PROC.sercon_8_0_o2[3]\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmdet[3]_net_1\, D => N_1064, Y => N_134);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_3_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        N_161_2, Y => N_161);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \un1_PCLK_count1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \un1_PCLK_count1_0_sqmuxa\, C => \PCLK_count1[1]_net_1\, 
        Y => CO1);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"FE0E")

      port map(A => \sercon_8_0_2[3]\, B => N_161, C => 
        un5_penable, D => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \sercon_9[3]\);
    
    PCLK_count1_0_sqmuxa_4 : CFG4
      generic map(INIT => x"0004")

      port map(A => \sercon[7]_net_1\, B => CO2_0, C => 
        \sercon[1]_net_1\, D => \sercon[0]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => \fsmsta[18]_net_1\, B => N_2177, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.CO2\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2_0);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2171, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    PCLK_count1_ov_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \PCLK_count1_ov_1_sqmuxa_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNIRHU61 : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        \pedetect\, C => un136_framesync, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \sercon[6]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_3_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \COREI2C_0_3_INT[0]\, B => N_2192, C => 
        \adrcomp_2_sqmuxa_i_0_0_0\, D => N_152, Y => 
        adrcomp_2_sqmuxa_i_0_2);
    
    \un2_framesync_1_1.CO1\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp_2_sqmuxa_i_a3_2\, B => 
        \framesync[1]_net_1\, Y => CO1_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"10")

      port map(A => fsmsta_8_23_351_i_0_1, B => N_2181, C => 
        N_1656, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        \serdat[0]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_9_509_0_1);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0D0F")

      port map(A => un92_fsmsta, B => \bsd7\, C => bsd7_9_iv_2, D
         => \un1_bsd7_1_sqmuxa[0]_net_1\, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \indelay[1]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \serdat_RNID9DU[4]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[4]_net_1\, B => \sercon[4]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[4]\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.ANC2\ : CFG3
      generic map(INIT => x"15")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => ANC2);
    
    \serSTA_WRITE_PROC.sersta_32_5[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[24]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_5[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_2177, B => N_172, Y => N_154);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    adrcomp_2_sqmuxa_i_a3 : CFG4
      generic map(INIT => x"D000")

      port map(A => mst, B => \fsmsta[23]_net_1\, C => N_2187, D
         => \adrcomp_2_sqmuxa_i_a3_3\, Y => N_152);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_0, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"4577")

      port map(A => \fsmsta[11]_net_1\, B => N_2177, C => N_2186, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[12]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    adrcomp_2_sqmuxa_i_0_0_0 : CFG2
      generic map(INIT => x"E")

      port map(A => un16_fsmmod, B => N_1586_1, Y => 
        \adrcomp_2_sqmuxa_i_0_0_0\);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2177, B => N_2178, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_3_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \fsmmod_ns_0_a4_0_1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \starto_en\, B => N_64, C => N_1040, D => 
        un115_fsmdet, Y => N_1059_1);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    adrcomp_2_sqmuxa_i_a3_2 : CFG2
      generic map(INIT => x"8")

      port map(A => \framesync[0]_net_1\, B => \nedetect\, Y => 
        \adrcomp_2_sqmuxa_i_a3_2\);
    
    un1_fsmsta_1_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => 
        \fsmsta[12]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => N_1470, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[14]_net_1\, 
        C => \fsmsta[18]_net_1\, Y => N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[0]\ : CFG4
      generic map(INIT => x"66F0")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync_7_m2[3]\, D => framesync_7_e2, Y => 
        \framesync_7[0]\);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    \sersta_RNI2S942[4]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        seradr0apb(7), Y => N_1221);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \un1_fsmsta_6\, B => un136_framesync, C => 
        \fsmsta_nxt_9_m_0[26]\, D => fsmsta_nxt_1_sqmuxa_18_s5_1, 
        Y => \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_1\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[2]_net_1\, C
         => un1_fsmmod, D => \fsmmod[0]_net_1\, Y => 
        SDAO_int_7_0_275_a5_1);
    
    \CLK_COUNTER1_PROC.un1_bclke_1.CO2\ : CFG3
      generic map(INIT => x"01")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[21]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_3_601_0_1, D => N_1717, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_ns_0_a4[5]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => \pedetect\, B => \SCLSCL\, C => un115_fsmdet, 
        D => \fsmmod[1]_net_1\, Y => N_1058);
    
    \fsmmod_ns_0_a4[0]\ : CFG4
      generic map(INIT => x"AAA2")

      port map(A => \fsmmod[6]_net_1\, B => \starto_en\, C => 
        N_1040, D => N_64, Y => N_1048);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    PCLKint_ff_RNIIH7R : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \serCON_WRITE_PROC.un3_penable\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_40, B => un3_penable_1, Y => un3_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_m2\ : CFG4
      generic map(INIT => x"C5C0")

      port map(A => \fsmsta[23]_net_1\, B => \fsmsta[9]_net_1\, C
         => N_2177, D => un1_fsmmod, Y => N_121);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \COREI2C_0_3_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_155, B => fsmsta_8_28_307_a3_0_0, C => 
        N_133, D => N_2181, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \sersta_32_i_a2_7[3]\, D => \COREI2C_0_3_INT[0]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    un1_fsmsta_1_i_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        Y => \un1_fsmsta_1_i_0_o2_0\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"00D0")

      port map(A => \PCLK_count1_ov_1_sqmuxa_1\, B => bclke, C
         => PCLK_count2_ov_6_1, D => \un1_PCLK_count1_0_sqmuxa\, 
        Y => \PCLK_count1_1_sqmuxa\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    serdat_2_sqmuxa : CFG4
      generic map(INIT => x"0020")

      port map(A => un92_fsmsta, B => un105_ens1, C => \pedetect\, 
        D => \COREI2C_0_3_INT[0]\, Y => \serdat_2_sqmuxa\);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_3_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        PCLK_count2_ov_6_1, C => CO1, D => \PCLK_count1_1_sqmuxa\, 
        Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => \fsmsta[16]_net_1\, B => N_2177, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_2177, B => \ack\, Y => N_155);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \sersta_RNIIB942[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => N_2186, B => N_2177, C => un136_framesync, D
         => N_82, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \sersta_32_4[1]\, B => m7_4, C => 
        \sersta_32_5[1]\, D => m7_5, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => un105_ens1_1, B => un3_penable, C => \ack\, D
         => CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \fsmsync_ns_i_o3_0_i_o2[5]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_64, B => \fsmsync[5]_net_1\, Y => N_68);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \un1_fsmsta_6\, B => un136_framesync, C => 
        \fsmsta_nxt_9_m_0[27]\, D => fsmsta_nxt_1_sqmuxa_24_s4_1, 
        Y => \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        \serdat[3]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[3]\ : CFG3
      generic map(INIT => x"6C")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[3]_net_1\, C => CO1_0, Y => 
        \framesync_7_enl_bm[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG3
      generic map(INIT => x"32")

      port map(A => fsmsta_8_5_555_a3_0_2, B => N_2181, C => 
        fsmsta_8_5_555_a3_2, Y => N_1665);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_3_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_3_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"3F20")

      port map(A => seradr0apb(0), B => \ack\, C => 
        un13_adrcompen, D => \adrcomp_2_sqmuxa_i_a2_1_5\, Y => 
        N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_3_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7[0]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_m2[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => N_1470);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \fsmsta_RNO[19]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_2199, B => un136_framesync, C => N_157, Y
         => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \COREI2C_0_3_INT[0]\, B => \sercon[5]_net_1\, 
        C => N_1041, D => \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => 
        N_1054);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        \serdat[5]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[6]\);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_0_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[4]_net_1\, Y => fsmsta_8_9_509_a4_0);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \fsmsta[14]_net_1\, D => \fsmsta[12]_net_1\, Y => 
        un25_fsmsta_1);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFDC")

      port map(A => N_2177, B => un16_fsmmod, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_3_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"3ACA")

      port map(A => \fsmdet[3]_net_1\, B => \framesync[1]_net_1\, 
        C => framesync_7_e2, D => \adrcomp_2_sqmuxa_i_a3_2\, Y
         => \framesync_7[1]\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => un16_fsmmod, B => \sercon_8_2[4]\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), D => un5_penable, Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => N_76, D => \fsmsync[4]_net_1\, Y => N_55_i_0);
    
    \serdat_RNI6UT91[6]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(6), B => \serdat[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => un91_ens1, B => N_2181, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \un1_PCLK_count1_0_sqmuxa\, D
         => \PCLK_count1_1_sqmuxa\, Y => \PCLK_count1_10[0]\);
    
    \serSTA_WRITE_PROC.sersta_32_4[0]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => \COREI2C_0_3_INT[0]\, B => N_127, C => 
        \fsmsta[9]_net_1\, Y => \sersta_32_4[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, Y => 
        un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    un1_PCLK_count1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"FF40")

      port map(A => \PCLK_count1[3]_net_1\, B => CO2, C => bclke, 
        D => \PCLK_count1_0_sqmuxa_3\, Y => 
        \un1_PCLK_count1_0_sqmuxa_1\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => mst, B => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"3AFF")

      port map(A => \COREI2C_0_3_SDAO[0]\, B => 
        \fsmsta[20]_net_1\, C => N_2177, D => N_2178, Y => 
        fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => \fsmmod[2]_net_1\, B => N_1064, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG3
      generic map(INIT => x"80")

      port map(A => un3_penable_1, B => un5_penable_1, C => N_40, 
        Y => un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    un1_PCLK_count1_0_sqmuxa_1_0 : CFG4
      generic map(INIT => x"080C")

      port map(A => \sercon[0]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => CO2, D => ANC2, Y => 
        \un1_PCLK_count1_0_sqmuxa_1_0\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG3
      generic map(INIT => x"20")

      port map(A => un137_framesync, B => \ack\, C => 
        un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_3_INT[0]\, 
        C => \sercon[5]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        \serdat[2]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => PCLK_count2_ov_6_0_a2_1_3, B => un16_fsmmod, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        \serdat[6]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[7]\);
    
    un1_counter_rst_3 : CFG2
      generic map(INIT => x"B")

      port map(A => \PCLK_count1_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, Y => \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_3_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"CACC")

      port map(A => \COREI2C_0_3_SDAO[0]\, B => 
        \fsmsta[13]_net_1\, C => N_2177, D => N_2196, Y => N_82);
    
    \fsmsta_RNO[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1656, B => N_2186, C => N_2181, D => N_124, 
        Y => N_1774_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_3_SDAO[0]\, Y => 
        N_172);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_4, B => N_145_2, C => 
        N_2177, D => fsmsta_8_20_379_i_0_a3_5, Y => N_145);
    
    adrcomp : SLE
      port map(D => N_2176_i_0, CLK => FAB_CCC_GL0, EN => 
        adrcomp_2_sqmuxa_i_0_2, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[19]_net_1\, 
        C => \fsmsta[4]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_4);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \fsmmod[0]_net_1\, B => \fsmdet[3]_net_1\, C
         => \fsmdet[1]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        N_1717);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_5\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => un135_ens1_2, Y => un135_ens1_5);
    
    \serCON_WRITE_PROC.un91_ens1_0_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \pedetect\, Y => un91_ens1);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[9]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    SDAO_int_RNI0N56 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_3_SDAO[0]\, Y => 
        COREI2C_0_3_SDAO_i(0));
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \PCLKint\, B => \PCLKint_ff\, C => N_1586_1, 
        D => \fsmmod[2]_net_1\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG3
      generic map(INIT => x"BF")

      port map(A => N_997, B => un70_fsmsta, C => 
        \fsmmod[4]_net_1\, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \fsmsync_RNO_0[1]\ : CFG4
      generic map(INIT => x"2232")

      port map(A => \fsmsync[2]_net_1\, B => N_997, C => 
        un70_fsmsta, D => N_68, Y => N_976_i_1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[26]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, Y
         => N_145_2);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => N_1665, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_68, B => \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \fsmmod[5]_net_1\, B => \nedetect\, C => 
        un115_fsmdet, D => N_1051, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_3_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    mst_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, Y
         => mst);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => un135_ens1_2, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_2181, B => fsmsta_8_2_647_i_0_0, C => 
        N_1656, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[20]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    un1_PCLK_count1_0_sqmuxa : CFG4
      generic map(INIT => x"EEEF")

      port map(A => \un1_PCLK_count1_0_sqmuxa_1\, B => 
        \un1_PCLK_count1_0_sqmuxa_0\, C => \sercon[7]_net_1\, D
         => \un1_PCLK_count1_0_sqmuxa_1_0\, Y => 
        \un1_PCLK_count1_0_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[22]\, B => un136_framesync, C
         => \fsmsta[22]_net_1\, D => N_2177, Y => \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_2, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \sersta_RNIUN942[3]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        \sercon[6]_net_1\, Y => N_1220);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_counter_rst_3\, D => 
        \un1_PCLK_count1_0_sqmuxa\, Y => \PCLK_count1_10[1]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_4\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, Y => un135_ens1_4);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG3
      generic map(INIT => x"F4")

      port map(A => \fsmmod[1]_net_1\, B => N_117_1, C => N_64, Y
         => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SCLInt\, B => \COREI2C_0_3_INT[0]\, C => 
        \bsd7_tmp\, Y => bsd7_tmp_i_m_1);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"FFEA")

      port map(A => un105_ens1, B => \serdat_2_sqmuxa\, C => 
        \sercon[6]_net_1\, D => \serdat_1_sqmuxa_1\, Y => 
        un1_serdat_2_sqmuxa_2);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \COREI2C_0_3_INT[0]\, B => N_1002, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_3_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_3_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"DCCC")

      port map(A => un105_ens1, B => \serdat_2_sqmuxa\, C => 
        \pedetect\, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_26_328_a3_0_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => \fsmsta[23]_net_1\, B => \adrcomp\, Y => N_26);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \serdat_RNIJFDU[7]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[7]_net_1\, B => \sercon[7]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \fsmdet[1]_net_1\, B => fsmsta_8_3_601_a4_0, 
        C => N_1656, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, C => 
        N_2193, D => N_172, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmmod[4]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, Y => N_1002);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_2\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => \fsmdet[3]_net_1\, B => \PWDATA_i_m_1[7]\, C
         => un105_ens1, D => bsd7_9_iv_1, Y => bsd7_9_iv_2);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_2_RNO\ : CFG4
      generic map(INIT => x"0002")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => \fsmdet[3]_net_1\, 
        D => \COREI2C_0_3_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[27]_net_1\, C => N_172, 
        Y => fsmsta_nxt_1_sqmuxa_24_s4_1);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[3]_net_1\, B => \serdat[2]_net_1\, C
         => \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[11]_net_1\, C
         => \fsmsta[7]_net_1\, D => \fsmsta[23]_net_1\, Y => m7_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[26]_net_1\, C => N_172, 
        Y => fsmsta_nxt_1_sqmuxa_18_s5_1);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        \serdat[4]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ack\, B => \adrcompen\, C => N_2177, D => 
        N_26, Y => fsmsta_8_5_555_a3_0_2);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_3_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3430")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1586_1, D => un1_fsmmod, Y => N_1624);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_3_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    un7_fsmsta_i_0_o2_RNIJDSC : CFG2
      generic map(INIT => x"1")

      port map(A => un57_fsmsta_1_0, B => N_2178, Y => N_191);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => \nedetect\, B => \COREI2C_0_3_INT[0]\, C => 
        \serdat[7]_net_1\, Y => \serdat_i_m_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_0_3\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[10]_net_1\, Y => fsmsta_8_3_601_a4_0);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    serdat_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \pedetect\, B => \sercon[6]_net_1\, C => 
        \un1_serdat40\, Y => \serdat_1_sqmuxa_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_1046, B => \fsmmod_ns_i_0[2]_net_1\, C => 
        N_1054, D => un115_fsmdet, Y => N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \CLK_COUNTER1_PROC.un12_pclk_count1_1.CO3\ : CFG4
      generic map(INIT => x"777F")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => un12_pclk_count1);
    
    adrcomp_RNO : CFG3
      generic map(INIT => x"15")

      port map(A => \adrcomp_2_sqmuxa_i_0_0_0\, B => 
        \COREI2C_0_3_INT[0]\, C => N_2192, Y => N_2176_i_0);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_am\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => un57_fsmsta, B => un105_ens1, C => \bsd7_tmp\, 
        D => bsd7_tmp_6_sn_m6_0, Y => bsd7_tmp_6_am_0);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_1[3]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_2179, B => \sercon[6]_net_1\, C => 
        un91_ens1, D => N_163, Y => \sercon_8_0_1[3]\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[23]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_5);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_3_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(2), B => seradr0apb(1), C => 
        \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => N_1449, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_3_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[16]_net_1\, 
        C => \fsmsta[20]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_2181, B => N_145, C => 
        fsmsta_8_20_379_i_0_o2_0, D => N_166, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_sm0, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[15]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[6]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \FSMSTA_SYNC_PROC.un137_framesync\ : CFG4
      generic map(INIT => x"0200")

      port map(A => un91_ens1, B => N_2181, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => un137_framesync);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_9_509_0_1, D => N_1717, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_126, B => N_80, C => un136_framesync, Y => 
        N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => un92_fsmsta, B => un105_ens1, C => 
        \serdat_i_m_1[7]\, D => bsd7_tmp_i_m_1, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \PCLKint\, B => \un151_framesync\, C => 
        \PCLKint_ff\, Y => \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \fsmdet[1]_net_1\, B => fsmsta_8_9_509_a4_0, 
        C => N_1656, D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"5444")

      port map(A => un115_fsmdet, B => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, C => \fsmmod[3]_net_1\, D
         => N_1034, Y => \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FDFF")

      port map(A => m7_4, B => \sersta_32_3[0]\, C => 
        \sersta_32_4[0]\, D => m7_5, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un135_ens1_4, B => un135_ens1_5, C => 
        \un1_fsmsta_1_i_0_o2_0\, D => un135_ens1_3, Y => 
        un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_2, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0501")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[6]_net_1\, C
         => \fsmmod[0]_net_1\, D => \adrcomp\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3[19]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => \SDAInt\, B => N_2178, C => N_2177, D => 
        N_191, Y => N_157);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG3
      generic map(INIT => x"80")

      port map(A => un3_penable_1, B => un105_ens1_1, C => N_40, 
        Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    \fsmsync_ns_i_a3_1_0_a2_2[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[3]_net_1\, C
         => \fsmmod[1]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_3_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_3\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[3]_net_1\, B => seradr0apb(4), Y => 
        un26_adrcompen_3);
    
    \sercon_RNIFBDU[5]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[5]_net_1\, B => \sercon[5]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    \fsmsync_RNO[1]\ : CFG4
      generic map(INIT => x"0D08")

      port map(A => \fsmsync[1]_net_1\, B => \SDAInt\, C => 
        N_1002, D => N_976_i_1, Y => N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1058, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_3_INT[0]\, 
        C => \fsmsta[28]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \sersta_RNIQJ942[2]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        seradr0apb(5), Y => N_1219);
    
    \serCON_WRITE_PROC.sercon_8_0_2[3]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \sercon[6]_net_1\, B => \COREI2C_0_3_INT[0]\, 
        C => \sercon_8_0_1[3]\, D => N_134, Y => 
        \sercon_8_0_2[3]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_3_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[3]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_enl_am[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG4
      generic map(INIT => x"ACCC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        \serdat[1]_net_1\, C => un3_penable, D => un105_ens1_1, Y
         => \serdat_9[2]\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[5]_net_1\, B => \fsmsync[2]_net_1\, 
        C => \fsmsync[1]_net_1\, D => \fsmsync[6]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => \nedetect\, B => N_117_1, C => 
        \fsmmod[4]_net_1\, Y => \fsmmod_ns_i_0[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_1586_1, B => N_2177, C => \fsmsta[8]_net_1\, 
        D => N_172, Y => fsmsta_8_5_555_a3_2);
    
    \fsmmod_ns_i_o3_0_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_3_INT[0]\, B => \sercon[4]_net_1\, 
        Y => N_997);
    
    adrcomp_2_sqmuxa_i_a3_2_0 : CFG3
      generic map(INIT => x"80")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \adrcomp_2_sqmuxa_i_a3_2\, Y
         => \adrcomp_2_sqmuxa_i_a3_2_0\);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG3
      generic map(INIT => x"02")

      port map(A => un137_framesync, B => \ack\, C => 
        un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_2);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_2 is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          COREI2C_0_3_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          un3_penable                  : in    std_logic;
          N_1217                       : out   std_logic;
          N_1218                       : out   std_logic;
          N_1220                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1221                       : out   std_logic;
          BIBUF_COREI2C_0_3_SDA_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_3_SCL_IO_Y   : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          bclke                        : in    std_logic;
          N_40                         : in    std_logic;
          un3_penable_1                : in    std_logic;
          un105_ens1_1                 : in    std_logic;
          un5_penable_1                : in    std_logic
        );

end COREI2C_2;

architecture DEF_ARCH of COREI2C_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_2
    port( COREI2C_0_3_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          seradr0apb                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          N_1217                       : out   std_logic;
          N_1218                       : out   std_logic;
          N_1220                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1221                       : out   std_logic;
          BIBUF_COREI2C_0_3_SDA_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_3_SCL_IO_Y   : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          bclke                        : in    std_logic := 'U';
          N_40                         : in    std_logic := 'U';
          un3_penable_1                : in    std_logic := 'U';
          un105_ens1_1                 : in    std_logic := 'U';
          un5_penable_1                : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_2
	Use entity work.COREI2CREAL_6_2(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_2
      port map(COREI2C_0_3_SDAO_i(0) => COREI2C_0_3_SDAO_i(0), 
        COREI2C_0_3_SCLO_i(0) => COREI2C_0_3_SCLO_i(0), 
        COREI2C_0_3_INT(0) => COREI2C_0_3_INT(0), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, N_1217 => N_1217, N_1218 => 
        N_1218, N_1220 => N_1220, N_1219 => N_1219, N_1221 => 
        N_1221, BIBUF_COREI2C_0_3_SDA_IO_Y => 
        BIBUF_COREI2C_0_3_SDA_IO_Y, BIBUF_COREI2C_0_3_SCL_IO_Y
         => BIBUF_COREI2C_0_3_SCL_IO_Y, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, bclke => bclke, N_40 => 
        N_40, un3_penable_1 => un3_penable_1, un105_ens1_1 => 
        un105_ens1_1, un5_penable_1 => un5_penable_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAPB3_MUXPTOB3 is

    port( GPOUT_reg                                   : in    std_logic_vector(31 downto 20);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 8);
          INTR_reg_m_0                                : in    std_logic;
          INTR_reg_m_9                                : in    std_logic;
          INTR_reg_m_4                                : in    std_logic;
          INTR_reg_m_7                                : in    std_logic;
          INTR_reg_m_1                                : in    std_logic;
          CoreAPB3_0_APBmslave7_PSELx                 : in    std_logic;
          N_440                                       : in    std_logic;
          un30_psel                                   : in    std_logic;
          N_438                                       : in    std_logic;
          N_439                                       : in    std_logic;
          N_435                                       : in    std_logic;
          N_441                                       : in    std_logic;
          N_437                                       : in    std_logic;
          N_436                                       : in    std_logic;
          N_338                                       : in    std_logic;
          N_333                                       : in    std_logic;
          N_310                                       : in    std_logic;
          N_419_mux                                   : in    std_logic;
          un3_prdata_o                                : in    std_logic;
          N_302                                       : in    std_logic;
          N_426_mux                                   : in    std_logic;
          N_345                                       : in    std_logic;
          N_421_mux                                   : in    std_logic;
          N_312                                       : in    std_logic;
          N_343                                       : in    std_logic;
          N_324                                       : in    std_logic;
          N_319                                       : in    std_logic;
          N_353                                       : in    std_logic;
          N_358                                       : in    std_logic;
          N_328                                       : in    std_logic
        );

end COREAPB3_MUXPTOB3;

architecture DEF_ARCH of COREAPB3_MUXPTOB3 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \PRDATA[17]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_333, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17));
    
    \PRDATA[30]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(30), C => N_439, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30));
    
    \PRDATA[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_338, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18));
    
    \PRDATA[8]\ : CFG4
      generic map(INIT => x"808C")

      port map(A => N_426_mux, B => CoreAPB3_0_APBmslave7_PSELx, 
        C => un3_prdata_o, D => N_345, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8));
    
    \PRDATA[31]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(31), C => INTR_reg_m_9, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31));
    
    \PRDATA[25]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(25), C => N_435, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25));
    
    \PRDATA[26]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(26), C => INTR_reg_m_4, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26));
    
    \PRDATA[24]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(24), C => N_436, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \PRDATA[20]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(20), C => N_438, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20));
    
    \PRDATA[29]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(29), C => INTR_reg_m_7, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29));
    
    \PRDATA[21]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(21), C => N_437, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21));
    
    \PRDATA[13]\ : CFG4
      generic map(INIT => x"808C")

      port map(A => N_421_mux, B => CoreAPB3_0_APBmslave7_PSELx, 
        C => un3_prdata_o, D => N_312, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13));
    
    \PRDATA[27]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(27), C => N_441, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27));
    
    \PRDATA[28]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(28), C => N_440, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28));
    
    \PRDATA[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_310, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12));
    
    \PRDATA[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_353, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9));
    
    \PRDATA[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_324, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \PRDATA[23]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(23), C => INTR_reg_m_1, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23));
    
    \PRDATA[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_328, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16));
    
    \PRDATA[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_319, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14));
    
    \PRDATA[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_358, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10));
    
    \PRDATA[19]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_343, B => CoreAPB3_0_APBmslave7_PSELx, Y
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19));
    
    \PRDATA[11]\ : CFG4
      generic map(INIT => x"808C")

      port map(A => N_419_mux, B => CoreAPB3_0_APBmslave7_PSELx, 
        C => un3_prdata_o, D => N_302, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11));
    
    \PRDATA[22]\ : CFG4
      generic map(INIT => x"A8A0")

      port map(A => CoreAPB3_0_APBmslave7_PSELx, B => 
        GPOUT_reg(22), C => INTR_reg_m_0, D => un30_psel, Y => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAPB3 is

    port( M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR  : in    std_logic_vector(15 downto 12);
          GPOUT_reg                                   : in    std_logic_vector(31 downto 20);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 8);
          CoreAPB3_0_APBmslave0_PADDR_8               : in    std_logic;
          CoreAPB3_0_APBmslave0_PADDR_7               : in    std_logic;
          CoreAPB3_0_APBmslave0_PADDR_0               : in    std_logic;
          CoreAPB3_0_APBmslave0_PADDR_6               : in    std_logic;
          CoreAPB3_0_APBmslave0_PADDR_5               : in    std_logic;
          INTR_reg_m_0                                : in    std_logic;
          INTR_reg_m_9                                : in    std_logic;
          INTR_reg_m_4                                : in    std_logic;
          INTR_reg_m_7                                : in    std_logic;
          INTR_reg_m_1                                : in    std_logic;
          N_8_0                                       : out   std_logic;
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : in    std_logic;
          m7_x                                        : out   std_logic;
          m46_1                                       : out   std_logic;
          N_122_i_1                                   : in    std_logic;
          N_122_i_0                                   : out   std_logic;
          N_92_i_1_1                                  : in    std_logic;
          N_92_i_0                                    : out   std_logic;
          N_48                                        : out   std_logic;
          m62_s                                       : in    std_logic;
          CONFIG_regror_28                            : in    std_logic;
          CONFIG_regror_29                            : in    std_logic;
          un561_psel_4                                : in    std_logic;
          N_1214                                      : in    std_logic;
          N_1215                                      : in    std_logic;
          N_1221                                      : in    std_logic;
          N_1219                                      : in    std_logic;
          N_1220                                      : in    std_logic;
          N_1218                                      : in    std_logic;
          N_1218_0                                    : in    std_logic;
          N_1218_1                                    : in    std_logic;
          N_1218_2                                    : in    std_logic;
          N_1216                                      : in    std_logic;
          N_1216_0                                    : in    std_logic;
          N_1216_1                                    : in    std_logic;
          N_1216_2                                    : in    std_logic;
          N_1216_3                                    : in    std_logic;
          N_1216_4                                    : in    std_logic;
          N_1214_0                                    : in    std_logic;
          N_1214_1                                    : in    std_logic;
          N_1214_2                                    : in    std_logic;
          N_1214_3                                    : in    std_logic;
          N_1214_4                                    : in    std_logic;
          N_1214_5                                    : in    std_logic;
          N_1217                                      : in    std_logic;
          N_1217_0                                    : in    std_logic;
          m71_1                                       : out   std_logic;
          N_1221_0                                    : in    std_logic;
          N_1221_1                                    : in    std_logic;
          N_1221_2                                    : in    std_logic;
          N_1221_3                                    : in    std_logic;
          N_1221_4                                    : in    std_logic;
          N_1221_5                                    : in    std_logic;
          N_1220_0                                    : in    std_logic;
          N_1220_1                                    : in    std_logic;
          N_1219_0                                    : in    std_logic;
          N_1219_1                                    : in    std_logic;
          N_1219_2                                    : in    std_logic;
          N_1219_3                                    : in    std_logic;
          N_1219_4                                    : in    std_logic;
          N_1219_5                                    : in    std_logic;
          N_1220_2                                    : in    std_logic;
          N_1220_3                                    : in    std_logic;
          N_1220_4                                    : in    std_logic;
          N_1220_5                                    : in    std_logic;
          N_1218_3                                    : in    std_logic;
          N_1218_4                                    : in    std_logic;
          N_1215_0                                    : in    std_logic;
          N_1215_1                                    : in    std_logic;
          N_1215_2                                    : in    std_logic;
          N_1215_3                                    : in    std_logic;
          N_1215_4                                    : in    std_logic;
          N_1215_5                                    : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE               : in    std_logic;
          CONFIG_rega23_1                             : in    std_logic;
          CoreAPB3_0_APBmslave7_PSELx                 : out   std_logic;
          N_1218_5                                    : in    std_logic;
          N_40                                        : out   std_logic;
          N_138                                       : out   std_logic;
          N_1216_5                                    : in    std_logic;
          N_43                                        : out   std_logic;
          un3_penable                                 : out   std_logic;
          un3_penable_0                               : out   std_logic;
          un3_penable_1                               : out   std_logic;
          un3_penable_2                               : out   std_logic;
          un3_penable_3                               : out   std_logic;
          un3_penable_4                               : out   std_logic;
          un3_penable_5                               : out   std_logic;
          N_24_0                                      : in    std_logic;
          N_137_i_0                                   : out   std_logic;
          N_37                                        : in    std_logic;
          N_107_i_0                                   : out   std_logic;
          N_53                                        : in    std_logic;
          N_62_i_0                                    : out   std_logic;
          N_58_0                                      : in    std_logic;
          N_38_i_0                                    : out   std_logic;
          N_63                                        : in    std_logic;
          N_23_0_i_0                                  : out   std_logic;
          N_440                                       : in    std_logic;
          un30_psel                                   : in    std_logic;
          N_438                                       : in    std_logic;
          N_439                                       : in    std_logic;
          N_435                                       : in    std_logic;
          N_441                                       : in    std_logic;
          N_437                                       : in    std_logic;
          N_436                                       : in    std_logic;
          N_338                                       : in    std_logic;
          N_333                                       : in    std_logic;
          N_310                                       : in    std_logic;
          N_419_mux                                   : in    std_logic;
          un3_prdata_o                                : in    std_logic;
          N_302                                       : in    std_logic;
          N_426_mux                                   : in    std_logic;
          N_345                                       : in    std_logic;
          N_421_mux                                   : in    std_logic;
          N_312                                       : in    std_logic;
          N_343                                       : in    std_logic;
          N_324                                       : in    std_logic;
          N_319                                       : in    std_logic;
          N_353                                       : in    std_logic;
          N_358                                       : in    std_logic;
          N_328                                       : in    std_logic
        );

end CoreAPB3;

architecture DEF_ARCH of CoreAPB3 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component COREAPB3_MUXPTOB3
    port( GPOUT_reg                                   : in    std_logic_vector(31 downto 20) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 8);
          INTR_reg_m_0                                : in    std_logic := 'U';
          INTR_reg_m_9                                : in    std_logic := 'U';
          INTR_reg_m_4                                : in    std_logic := 'U';
          INTR_reg_m_7                                : in    std_logic := 'U';
          INTR_reg_m_1                                : in    std_logic := 'U';
          CoreAPB3_0_APBmslave7_PSELx                 : in    std_logic := 'U';
          N_440                                       : in    std_logic := 'U';
          un30_psel                                   : in    std_logic := 'U';
          N_438                                       : in    std_logic := 'U';
          N_439                                       : in    std_logic := 'U';
          N_435                                       : in    std_logic := 'U';
          N_441                                       : in    std_logic := 'U';
          N_437                                       : in    std_logic := 'U';
          N_436                                       : in    std_logic := 'U';
          N_338                                       : in    std_logic := 'U';
          N_333                                       : in    std_logic := 'U';
          N_310                                       : in    std_logic := 'U';
          N_419_mux                                   : in    std_logic := 'U';
          un3_prdata_o                                : in    std_logic := 'U';
          N_302                                       : in    std_logic := 'U';
          N_426_mux                                   : in    std_logic := 'U';
          N_345                                       : in    std_logic := 'U';
          N_421_mux                                   : in    std_logic := 'U';
          N_312                                       : in    std_logic := 'U';
          N_343                                       : in    std_logic := 'U';
          N_324                                       : in    std_logic := 'U';
          N_319                                       : in    std_logic := 'U';
          N_353                                       : in    std_logic := 'U';
          N_358                                       : in    std_logic := 'U';
          N_328                                       : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \m7_sx\, \m7_2_0\, \N_8_0\, \m83_bm\, m91_d_0_1, 
        \m83_am\, \m91_d_0\, N_88, N_87, N_53_0, \m61_d_0_1_0\, 
        N_50, \m61_d_0\, N_58, N_57, \m121_d\, m46_1_net_1, 
        N_92_i_1, \m61_s\, \N_48\, \m17_1\, \m22_d_1_1_1\, 
        \m22_d_1_1\, \m22_d_1_0\, \m22_d\, \m13_1\, \m22_d_1_0_1\, 
        \m10_1\, \m32_ns_1\, \m37_d_1_1_1\, \m37_d_1_1\, 
        \m37_d_1_0\, \m37_d\, \m28_ns_1\, \m37_d_1_0_1\, 
        \m25_ns_1\, \m131_1\, \m136_d_1_1_1\, \m136_d_1_1\, 
        \m136_d_1_0\, \m136_d\, \m127_1\, \m136_d_1_0_1\, 
        \m124_1\, \m101_1\, \m106_d_1_1_1\, \m106_d_1_1\, 
        \m106_d_1_0\, \m106_d\, \m97_ns_1\, \m106_d_1_0_1\, 
        \m94_ns_1\, \m116_1\, \m121_d_1_1_1\, \m121_d_1_1\, 
        \m121_d_1_0\, \m112_ns_1\, \m121_d_1_0_1\, \m109_ns_1\, 
        \m83_am_1\, \m83_bm_1\, \m49_1\, \m52_1\, \m56_1\, 
        \m86_ns_1\, \m7_2\, \m3_3\, \CoreAPB3_0_APBmslave7_PSELx\, 
        N_157_mux, GND_net_1, VCC_net_1 : std_logic;

    for all : COREAPB3_MUXPTOB3
	Use entity work.COREAPB3_MUXPTOB3(DEF_ARCH);
begin 

    N_8_0 <= \N_8_0\;
    m46_1 <= m46_1_net_1;
    N_48 <= \N_48\;
    CoreAPB3_0_APBmslave7_PSELx <= \CoreAPB3_0_APBmslave7_PSELx\;

    \iPSELS_raw_1_0_a2_0_RNIT2OO1[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \N_48\, B => un561_psel_4, C => \m3_3\, Y => 
        N_157_mux);
    
    m17_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1214_0, C => N_1214_1, Y => \m17_1\);
    
    m22_d_1_0_1 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        un561_psel_4, C => \N_8_0\, Y => \m22_d_1_0_1\);
    
    m7_sx : CFG3
      generic map(INIT => x"FD")

      port map(A => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, B
         => M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15), C => 
        CoreAPB3_0_APBmslave0_PADDR_7, Y => \m7_sx\);
    
    m106_d_1_0_1 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        un561_psel_4, C => \N_8_0\, Y => \m106_d_1_0_1\);
    
    m37_d_1_0 : CFG4
      generic map(INIT => x"4070")

      port map(A => \m28_ns_1\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        \m37_d_1_0_1\, D => \m25_ns_1\, Y => \m37_d_1_0\);
    
    m32_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1215_4, C => N_1215_5, Y => \m32_ns_1\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_2[0]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_5);
    
    \m71_1\ : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1217, C => N_1217_0, Y => m71_1);
    
    m121_d_1_1_1 : CFG4
      generic map(INIT => x"3010")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PADDR_0, C => un561_psel_4, D => 
        N_1220, Y => \m121_d_1_1_1\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_5[0]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_3);
    
    m57 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1216_5, B => \N_8_0\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_58);
    
    m124_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1221_0, C => N_1221_1, Y => \m124_1\);
    
    u_mux_p_to_b3 : COREAPB3_MUXPTOB3
      port map(GPOUT_reg(31) => GPOUT_reg(31), GPOUT_reg(30) => 
        GPOUT_reg(30), GPOUT_reg(29) => GPOUT_reg(29), 
        GPOUT_reg(28) => GPOUT_reg(28), GPOUT_reg(27) => 
        GPOUT_reg(27), GPOUT_reg(26) => GPOUT_reg(26), 
        GPOUT_reg(25) => GPOUT_reg(25), GPOUT_reg(24) => 
        GPOUT_reg(24), GPOUT_reg(23) => GPOUT_reg(23), 
        GPOUT_reg(22) => GPOUT_reg(22), GPOUT_reg(21) => 
        GPOUT_reg(21), GPOUT_reg(20) => GPOUT_reg(20), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        INTR_reg_m_0 => INTR_reg_m_0, INTR_reg_m_9 => 
        INTR_reg_m_9, INTR_reg_m_4 => INTR_reg_m_4, INTR_reg_m_7
         => INTR_reg_m_7, INTR_reg_m_1 => INTR_reg_m_1, 
        CoreAPB3_0_APBmslave7_PSELx => 
        \CoreAPB3_0_APBmslave7_PSELx\, N_440 => N_440, un30_psel
         => un30_psel, N_438 => N_438, N_439 => N_439, N_435 => 
        N_435, N_441 => N_441, N_437 => N_437, N_436 => N_436, 
        N_338 => N_338, N_333 => N_333, N_310 => N_310, N_419_mux
         => N_419_mux, un3_prdata_o => un3_prdata_o, N_302 => 
        N_302, N_426_mux => N_426_mux, N_345 => N_345, N_421_mux
         => N_421_mux, N_312 => N_312, N_343 => N_343, N_324 => 
        N_324, N_319 => N_319, N_353 => N_353, N_358 => N_358, 
        N_328 => N_328);
    
    m61_d_0 : CFG4
      generic map(INIT => x"F2C2")

      port map(A => N_53_0, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => 
        \m61_d_0_1_0\, D => N_50, Y => \m61_d_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    m97_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1219_4, C => N_1219_5, Y => \m97_ns_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIV3DT1_1[0]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \N_48\, B => \m7_2\, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        N_138);
    
    m83_am_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1218, C => N_1218_0, Y => \m83_am_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIJB8SN2[0]\ : CFG4
      generic map(INIT => x"1D11")

      port map(A => \m121_d\, B => m46_1_net_1, C => N_92_i_1, D
         => N_122_i_1, Y => N_122_i_0);
    
    m37_d_1_1_1 : CFG4
      generic map(INIT => x"3010")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PADDR_0, C => un561_psel_4, D => 
        N_1215, Y => \m37_d_1_1_1\);
    
    m83_bm_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1218_1, C => N_1218_2, Y => \m83_bm_1\);
    
    \m7_x\ : CFG3
      generic map(INIT => x"04")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_8, B => \m7_2_0\, 
        C => CoreAPB3_0_APBmslave0_PADDR_7, Y => m7_x);
    
    m49 : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m49_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_50);
    
    m22_d_1_1_1 : CFG4
      generic map(INIT => x"3010")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PADDR_0, C => un561_psel_4, D => 
        N_1214, Y => \m22_d_1_1_1\);
    
    m91_d_0 : CFG4
      generic map(INIT => x"F2C2")

      port map(A => \m83_bm\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => 
        m91_d_0_1, D => \m83_am\, Y => \m91_d_0\);
    
    m7_2 : CFG4
      generic map(INIT => x"0001")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_5, B => 
        CoreAPB3_0_APBmslave0_PADDR_7, C => 
        CoreAPB3_0_APBmslave0_PADDR_8, D => 
        CoreAPB3_0_APBmslave0_PADDR_6, Y => \m7_2\);
    
    m37_d_1_1 : CFG4
      generic map(INIT => x"73FF")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        \N_8_0\, C => \m32_ns_1\, D => \m37_d_1_1_1\, Y => 
        \m37_d_1_1\);
    
    m106_d_1_1_1 : CFG4
      generic map(INIT => x"3010")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PADDR_0, C => un561_psel_4, D => 
        N_1219, Y => \m106_d_1_1_1\);
    
    m136_d_1_0_1 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        un561_psel_4, C => \N_8_0\, Y => \m136_d_1_0_1\);
    
    \iPSELS_raw_1_0_a2_0[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, Y => \N_48\);
    
    m49_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1216, C => N_1216_0, Y => \m49_1\);
    
    m136_d : CFG3
      generic map(INIT => x"8D")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \m136_d_1_1\, C => \m136_d_1_0\, Y => \m136_d\);
    
    m131_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1221_4, C => N_1221_5, Y => \m131_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    m37_d : CFG3
      generic map(INIT => x"8D")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \m37_d_1_1\, C => \m37_d_1_0\, Y => \m37_d\);
    
    m28_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1215_2, C => N_1215_3, Y => \m28_ns_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIV3DT1[0]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \N_48\, B => \m7_2\, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => N_43);
    
    \iPSELS_raw_1_0_a2_0_RNIGMI01[0]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \N_48\, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        \CoreAPB3_0_APBmslave7_PSELx\);
    
    m112_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1220_4, C => N_1220_5, Y => \m112_ns_1\);
    
    m10_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1214_4, C => N_1214_5, Y => \m10_1\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2[0]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable);
    
    m86_ns : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m86_ns_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_87);
    
    m83_bm : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m83_bm_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        \m83_bm\);
    
    m3_3 : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        CoreAPB3_0_APBmslave0_PWRITE, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => CONFIG_rega23_1, Y
         => \m3_3\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_1[0]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_1);
    
    m7_2_0 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_6, B => 
        CoreAPB3_0_APBmslave0_PADDR_5, Y => \m7_2_0\);
    
    m127_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1221_2, C => N_1221_3, Y => \m127_1\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_0[0]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_0);
    
    \iPSELS_raw_1_0_a2_0_RNIQ6Q0S2[0]\ : CFG4
      generic map(INIT => x"3505")

      port map(A => \m91_d_0\, B => N_92_i_1, C => \m61_s\, D => 
        N_92_i_1_1, Y => N_92_i_0);
    
    m56_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1216_3, C => N_1216_4, Y => \m56_1\);
    
    m52_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1216_1, C => N_1216_2, Y => \m52_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIR108Q2[0]\ : CFG4
      generic map(INIT => x"038B")

      port map(A => \N_48\, B => m46_1_net_1, C => \m106_d\, D
         => N_37, Y => N_107_i_0);
    
    m136_d_1_0 : CFG4
      generic map(INIT => x"4070")

      port map(A => \m127_1\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        \m136_d_1_0_1\, D => \m124_1\, Y => \m136_d_1_0\);
    
    m106_d_1_0 : CFG4
      generic map(INIT => x"4070")

      port map(A => \m97_ns_1\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        \m106_d_1_0_1\, D => \m94_ns_1\, Y => \m106_d_1_0\);
    
    m22_d : CFG3
      generic map(INIT => x"8D")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \m22_d_1_1\, C => \m22_d_1_0\, Y => \m22_d\);
    
    \iPSELS_raw_1_0_a2_0_RNIV3DT1_0[0]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \N_48\, B => \m7_2\, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => N_40);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_4[0]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_2);
    
    m87 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1218_5, B => \N_8_0\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_88);
    
    m136_d_1_1_1 : CFG4
      generic map(INIT => x"3010")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PADDR_0, C => un561_psel_4, D => 
        N_1221, Y => \m136_d_1_1_1\);
    
    m91_d_0_1_0 : CFG4
      generic map(INIT => x"5D19")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => N_88, 
        D => N_87, Y => m91_d_0_1);
    
    \iPSELS_raw_1_0_a2_0_RNIR78AQ2[0]\ : CFG4
      generic map(INIT => x"038B")

      port map(A => \N_48\, B => m46_1_net_1, C => \m136_d\, D
         => N_24_0, Y => N_137_i_0);
    
    m83_am : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m83_am_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        \m83_am\);
    
    m116_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1220_0, C => N_1220_1, Y => \m116_1\);
    
    \iPSELS_raw_1_0_a2_0_RNI82BSB2[0]\ : CFG4
      generic map(INIT => x"038B")

      port map(A => \N_48\, B => m46_1_net_1, C => \m22_d\, D => 
        N_63, Y => N_23_0_i_0);
    
    m7 : CFG3
      generic map(INIT => x"10")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_8, B => \m7_sx\, 
        C => \m7_2_0\, Y => \N_8_0\);
    
    m13_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1214_2, C => N_1214_3, Y => \m13_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIH20GQ1[0]\ : CFG4
      generic map(INIT => x"555D")

      port map(A => \N_48\, B => m62_s, C => CONFIG_regror_28, D
         => CONFIG_regror_29, Y => N_92_i_1);
    
    m86_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1218_3, C => N_1218_4, Y => \m86_ns_1\);
    
    m121_d_1_0_1 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        un561_psel_4, C => \N_8_0\, Y => \m121_d_1_0_1\);
    
    \iPSELS_raw_1_0_a2_0_RNI1M53G2[0]\ : CFG4
      generic map(INIT => x"3505")

      port map(A => \m61_d_0\, B => N_53, C => \m61_s\, D => 
        \N_48\, Y => N_62_i_0);
    
    m106_d : CFG3
      generic map(INIT => x"8D")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \m106_d_1_1\, C => \m106_d_1_0\, Y => \m106_d\);
    
    m101_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1219_0, C => N_1219_1, Y => \m101_1\);
    
    m52 : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m52_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_53_0);
    
    \m46_1\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), Y => 
        m46_1_net_1);
    
    m37_d_1_0_1 : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR_0, B => 
        un561_psel_4, C => \N_8_0\, Y => \m37_d_1_0_1\);
    
    m22_d_1_1 : CFG4
      generic map(INIT => x"73FF")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        \N_8_0\, C => \m17_1\, D => \m22_d_1_1_1\, Y => 
        \m22_d_1_1\);
    
    m136_d_1_1 : CFG4
      generic map(INIT => x"73FF")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        \N_8_0\, C => \m131_1\, D => \m136_d_1_1_1\, Y => 
        \m136_d_1_1\);
    
    m94_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1219_2, C => N_1219_3, Y => \m94_ns_1\);
    
    m109_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1220_2, C => N_1220_3, Y => \m109_ns_1\);
    
    m106_d_1_1 : CFG4
      generic map(INIT => x"73FF")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        \N_8_0\, C => \m101_1\, D => \m106_d_1_1_1\, Y => 
        \m106_d_1_1\);
    
    m121_d_1_1 : CFG4
      generic map(INIT => x"73FF")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        \N_8_0\, C => \m116_1\, D => \m121_d_1_1_1\, Y => 
        \m121_d_1_1\);
    
    \iPSELS_raw_1_0_a2_0_RNIHBBSB2[0]\ : CFG4
      generic map(INIT => x"038B")

      port map(A => \N_48\, B => m46_1_net_1, C => \m37_d\, D => 
        N_58_0, Y => N_38_i_0);
    
    m61_s : CFG3
      generic map(INIT => x"80")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), Y => 
        \m61_s\);
    
    m22_d_1_0 : CFG4
      generic map(INIT => x"4070")

      port map(A => \m13_1\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        \m22_d_1_0_1\, D => \m10_1\, Y => \m22_d_1_0\);
    
    \iPSELS_raw_1_0_a2_0_RNICGIL2_3[0]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        N_157_mux, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un3_penable_4);
    
    m56 : CFG4
      generic map(INIT => x"FDFF")

      port map(A => \N_8_0\, B => \m56_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR_0, D => un561_psel_4, Y => 
        N_57);
    
    m121_d : CFG3
      generic map(INIT => x"8D")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        \m121_d_1_1\, C => \m121_d_1_0\, Y => \m121_d\);
    
    m61_d_0_1_0 : CFG4
      generic map(INIT => x"5D19")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), C => N_58, 
        D => N_57, Y => \m61_d_0_1_0\);
    
    m25_ns_1 : CFG3
      generic map(INIT => x"27")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), B => 
        N_1215_0, C => N_1215_1, Y => \m25_ns_1\);
    
    m121_d_1_0 : CFG4
      generic map(INIT => x"4070")

      port map(A => \m112_ns_1\, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), C => 
        \m121_d_1_0_1\, D => \m109_ns_1\, Y => \m121_d_1_0\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreGPIO is

    port( CoreAPB3_0_APBmslave0_PWDATA  : in    std_logic_vector(31 downto 0);
          GPIO_IN_c                     : in    std_logic_vector(19 downto 4);
          CoreAPB3_0_APBmslave0_PADDR   : in    std_logic_vector(7 downto 0);
          GPIO_OUT_c                    : out   std_logic_vector(2 downto 1);
          GPOUT_reg_3                   : out   std_logic;
          GPOUT_reg_31                  : out   std_logic;
          GPOUT_reg_30                  : out   std_logic;
          GPOUT_reg_29                  : out   std_logic;
          GPOUT_reg_28                  : out   std_logic;
          GPOUT_reg_27                  : out   std_logic;
          GPOUT_reg_26                  : out   std_logic;
          GPOUT_reg_25                  : out   std_logic;
          GPOUT_reg_24                  : out   std_logic;
          GPOUT_reg_23                  : out   std_logic;
          GPOUT_reg_22                  : out   std_logic;
          GPOUT_reg_21                  : out   std_logic;
          GPOUT_reg_20                  : out   std_logic;
          INTR_reg_m_0                  : out   std_logic;
          INTR_reg_m_9                  : out   std_logic;
          INTR_reg_m_4                  : out   std_logic;
          INTR_reg_m_7                  : out   std_logic;
          INTR_reg_m_1                  : out   std_logic;
          MSS_READY                     : in    std_logic;
          FAB_CCC_GL0                   : in    std_logic;
          un30_psel                     : out   std_logic;
          m62_s                         : out   std_logic;
          un3_prdata_o                  : out   std_logic;
          CONFIG_regror_29              : out   std_logic;
          CONFIG_regror_28              : out   std_logic;
          N_24_0                        : out   std_logic;
          N_53                          : out   std_logic;
          N_58                          : out   std_logic;
          N_37                          : out   std_logic;
          N_122_i_1                     : out   std_logic;
          N_63                          : out   std_logic;
          N_92_i_1_1                    : out   std_logic;
          N_47                          : out   std_logic;
          N_310                         : out   std_logic;
          N_333                         : out   std_logic;
          N_338                         : out   std_logic;
          N_343                         : out   std_logic;
          N_319                         : out   std_logic;
          N_6186                        : out   std_logic;
          N_324                         : out   std_logic;
          N_353                         : out   std_logic;
          N_358                         : out   std_logic;
          N_328                         : out   std_logic;
          N_419_mux                     : out   std_logic;
          N_426_mux                     : out   std_logic;
          USB_RST_c                     : out   std_logic;
          N_421_mux                     : out   std_logic;
          CONFIG_rega23_1               : out   std_logic;
          CONFIG_rega20_2               : in    std_logic;
          N_48_1                        : in    std_logic;
          m46_1_0                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE  : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE : in    std_logic;
          CoreAPB3_0_APBmslave7_PSELx   : in    std_logic;
          N_438                         : out   std_logic;
          N_440                         : out   std_logic;
          N_439                         : out   std_logic;
          N_435                         : out   std_logic;
          N_441                         : out   std_logic;
          N_437                         : out   std_logic;
          N_436                         : out   std_logic;
          N_302                         : out   std_logic;
          N_345                         : out   std_logic;
          N_312                         : out   std_logic
        );

end CoreGPIO;

architecture DEF_ARCH of CoreGPIO is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM64x18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_ADDR_CLK    : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ADDR_SRST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_ADDR_ARST_N : in    std_logic := 'U';
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_ADDR_EN     : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          B_ADDR_CLK    : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ADDR_SRST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_ADDR_ARST_N : in    std_logic := 'U';
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_ADDR_EN     : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_CLK         : in    std_logic := 'U';
          C_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          C_WEN         : in    std_logic := 'U';
          C_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_ADDR_LAT    : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_EN          : in    std_logic := 'U';
          B_ADDR_LAT    : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          C_EN          : in    std_logic := 'U';
          C_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \CONFIG_reg_28[7]_net_1\, VCC_net_1, un822_psel, 
        GND_net_1, \CONFIG_reg_14[7]_net_1\, un416_psel, 
        \CONFIG_reg_13[5]_net_1\, un387_psel, 
        \CONFIG_reg_13[6]_net_1\, \CONFIG_reg_13[7]_net_1\, 
        \CONFIG_reg_31[5]_net_1\, un909_psel, 
        \CONFIG_reg_31[6]_net_1\, \CONFIG_reg_31[7]_net_1\, 
        \CONFIG_reg_30[5]_net_1\, un880_psel, 
        \CONFIG_reg_30[6]_net_1\, \CONFIG_reg_30[7]_net_1\, 
        \CONFIG_reg_29[5]_net_1\, un851_psel, 
        \CONFIG_reg_29[6]_net_1\, \CONFIG_reg_29[7]_net_1\, 
        \CONFIG_reg_28[5]_net_1\, \CONFIG_reg_28[6]_net_1\, 
        \CONFIG_reg_19[7]_net_1\, un561_psel, 
        \CONFIG_reg_18[5]_net_1\, un532_psel, 
        \CONFIG_reg_18[6]_net_1\, \CONFIG_reg_18[7]_net_1\, 
        \CONFIG_reg_17[5]_net_1\, un503_psel, 
        \CONFIG_reg_17[6]_net_1\, \CONFIG_reg_17[7]_net_1\, 
        \CONFIG_reg_16[5]_net_1\, un474_psel, 
        \CONFIG_reg_16[6]_net_1\, \CONFIG_reg_16[7]_net_1\, 
        \CONFIG_reg_15[5]_net_1\, un445_psel, 
        \CONFIG_reg_15[6]_net_1\, \CONFIG_reg_15[7]_net_1\, 
        \CONFIG_reg_14[5]_net_1\, \CONFIG_reg_14[6]_net_1\, 
        \CONFIG_reg_24[7]_net_1\, un706_psel, 
        \CONFIG_reg_23[5]_net_1\, un677_psel, 
        \CONFIG_reg_23[6]_net_1\, \CONFIG_reg_23[7]_net_1\, 
        \CONFIG_reg_22[5]_net_1\, un648_psel, 
        \CONFIG_reg_22[6]_net_1\, \CONFIG_reg_22[7]_net_1\, 
        \CONFIG_reg_21[5]_net_1\, un619_psel, 
        \CONFIG_reg_21[6]_net_1\, \CONFIG_reg_21[7]_net_1\, 
        \CONFIG_reg_20[5]_net_1\, un590_psel, 
        \CONFIG_reg_20[6]_net_1\, \CONFIG_reg_20[7]_net_1\, 
        \CONFIG_reg_19[5]_net_1\, \CONFIG_reg_19[6]_net_1\, 
        \CONFIG_reg_0[7]_net_1\, un11_psel, 
        \CONFIG_reg_31[0]_net_1\, \CONFIG_reg_31[3]_net_1\, 
        \CONFIG_reg_30[3]_net_1\, \CONFIG_reg_27[5]_net_1\, 
        un793_psel, \CONFIG_reg_27[6]_net_1\, 
        \CONFIG_reg_27[7]_net_1\, \CONFIG_reg_26[5]_net_1\, 
        un764_psel, \CONFIG_reg_26[6]_net_1\, 
        \CONFIG_reg_26[7]_net_1\, \CONFIG_reg_25[5]_net_1\, 
        un735_psel, \CONFIG_reg_25[6]_net_1\, 
        \CONFIG_reg_25[7]_net_1\, \CONFIG_reg_24[5]_net_1\, 
        \CONFIG_reg_24[6]_net_1\, \CONFIG_reg_5[7]_net_1\, 
        un156_psel, \CONFIG_reg_4[5]_net_1\, un127_psel, 
        \CONFIG_reg_4[6]_net_1\, \CONFIG_reg_4[7]_net_1\, 
        \CONFIG_reg_3[5]_net_1\, un98_psel, 
        \CONFIG_reg_3[6]_net_1\, \CONFIG_reg_3[7]_net_1\, 
        \CONFIG_reg_2[5]_net_1\, un69_psel, 
        \CONFIG_reg_2[6]_net_1\, \CONFIG_reg_2[7]_net_1\, 
        \CONFIG_reg_1[5]_net_1\, un41_psel, 
        \CONFIG_reg_1[6]_net_1\, \CONFIG_reg_1[7]_net_1\, 
        \CONFIG_reg_0[5]_net_1\, \CONFIG_reg_0[6]_net_1\, 
        \CONFIG_reg_10[7]_net_1\, un300_psel, 
        \CONFIG_reg_9[5]_net_1\, un271_psel, 
        \CONFIG_reg_9[6]_net_1\, \CONFIG_reg_9[7]_net_1\, 
        \CONFIG_reg_8[5]_net_1\, un242_psel, 
        \CONFIG_reg_8[6]_net_1\, \CONFIG_reg_8[7]_net_1\, 
        \CONFIG_reg_7[5]_net_1\, un214_psel, 
        \CONFIG_reg_7[6]_net_1\, \CONFIG_reg_7[7]_net_1\, 
        \CONFIG_reg_6[5]_net_1\, un185_psel, 
        \CONFIG_reg_6[6]_net_1\, \CONFIG_reg_6[7]_net_1\, 
        \CONFIG_reg_5[5]_net_1\, \CONFIG_reg_5[6]_net_1\, 
        \CONFIG_reg_18[3]_net_1\, \CONFIG_reg_17[1]_net_1\, 
        \CONFIG_reg_17[3]_net_1\, \CONFIG_reg_16[1]_net_1\, 
        \CONFIG_reg_16[3]_net_1\, \CONFIG_reg_15[1]_net_1\, 
        \CONFIG_reg_15[3]_net_1\, \CONFIG_reg_12[5]_net_1\, 
        un358_psel, \CONFIG_reg_12[6]_net_1\, 
        \CONFIG_reg_12[7]_net_1\, \CONFIG_reg_11[5]_net_1\, 
        un329_psel, \CONFIG_reg_11[6]_net_1\, 
        \CONFIG_reg_11[7]_net_1\, \CONFIG_reg_10[5]_net_1\, 
        \CONFIG_reg_10[6]_net_1\, \CONFIG_reg_1[3]_net_1\, 
        \CONFIG_reg_0[3]_net_1\, \CONFIG_reg_29[3]_net_1\, 
        \CONFIG_reg_28[3]_net_1\, \CONFIG_reg_27[3]_net_1\, 
        \CONFIG_reg_26[3]_net_1\, \CONFIG_reg_25[3]_net_1\, 
        \CONFIG_reg_24[3]_net_1\, \CONFIG_reg_23[3]_net_1\, 
        \CONFIG_reg_22[3]_net_1\, \CONFIG_reg_21[3]_net_1\, 
        \CONFIG_reg_20[3]_net_1\, \CONFIG_reg_19[1]_net_1\, 
        \CONFIG_reg_19[3]_net_1\, \CONFIG_reg_18[1]_net_1\, 
        \CONFIG_reg_9[3]_net_1\, \CONFIG_reg_8[1]_net_1\, 
        \CONFIG_reg_8[3]_net_1\, \CONFIG_reg_7[1]_net_1\, 
        \CONFIG_reg_7[3]_net_1\, \CONFIG_reg_6[1]_net_1\, 
        \CONFIG_reg_6[3]_net_1\, \CONFIG_reg_5[1]_net_1\, 
        \CONFIG_reg_5[3]_net_1\, \CONFIG_reg_4[1]_net_1\, 
        \CONFIG_reg_4[3]_net_1\, \CONFIG_reg_3[3]_net_1\, 
        \CONFIG_reg_2[0]_net_1\, \CONFIG_reg_2[3]_net_1\, 
        \CONFIG_reg_1[0]_net_1\, \CONFIG_reg_14[1]_net_1\, 
        \CONFIG_reg_14[3]_net_1\, \CONFIG_reg_13[1]_net_1\, 
        \CONFIG_reg_13[3]_net_1\, \CONFIG_reg_12[1]_net_1\, 
        \CONFIG_reg_12[3]_net_1\, \CONFIG_reg_11[1]_net_1\, 
        \CONFIG_reg_11[3]_net_1\, \CONFIG_reg_10[1]_net_1\, 
        \CONFIG_reg_10[3]_net_1\, \CONFIG_reg_9[1]_net_1\, 
        CONFIG_regro_27, CONFIG_regro_28, CONFIG_regro_29, 
        CONFIG_regro_30, CONFIG_regro_31, CONFIG_regro_22, 
        CONFIG_regro_23, CONFIG_regro_24, CONFIG_regro_25, 
        CONFIG_regro_26, CONFIG_regro_17, CONFIG_regro_18, 
        CONFIG_regro_19, CONFIG_regro_20, CONFIG_regro_21, 
        CONFIG_regro_12, CONFIG_regro_13, CONFIG_regro_14, 
        CONFIG_regro_15, CONFIG_regro_16, CONFIG_regro_7, 
        CONFIG_regro_8, CONFIG_regro_9, CONFIG_regro_10, 
        CONFIG_regro_11, CONFIG_regro_2, CONFIG_regro_3, 
        CONFIG_regro_4, CONFIG_regro_5, CONFIG_regro_6, 
        CONFIG_regro_0, CONFIG_regro_1, \GPOUT_reg[4]_net_1\, 
        N_51_i_0, \GPOUT_reg[2]_net_1\, \GPOUT_reg[1]_net_1\, 
        \GPOUT_reg[0]_net_1\, \GPOUT_reg[19]_net_1\, 
        \GPOUT_reg[18]_net_1\, \GPOUT_reg[17]_net_1\, 
        \GPOUT_reg[16]_net_1\, \GPOUT_reg[15]_net_1\, 
        \GPOUT_reg[14]_net_1\, \GPOUT_reg[13]_net_1\, 
        \GPOUT_reg[12]_net_1\, \GPOUT_reg[11]_net_1\, 
        \GPOUT_reg[10]_net_1\, \GPOUT_reg[9]_net_1\, 
        \GPOUT_reg[8]_net_1\, \GPOUT_reg[7]_net_1\, 
        \GPOUT_reg[6]_net_1\, \GPOUT_reg[5]_net_1\, 
        \edge_pos[6]_net_1\, \edge_pos_67_iv_i_0[6]\, 
        edge_pos_2_sqmuxa_388_i_0, \edge_pos[5]_net_1\, 
        \edge_pos_57_iv_i_0[5]\, edge_pos_2_sqmuxa_389_i_0, 
        \edge_pos[4]_net_1\, \edge_pos_47_iv_i_0[4]\, 
        edge_pos_2_sqmuxa_375_i_0, \GPOUT_reg_31\, 
        \edge_neg[5]_net_1\, \edge_neg_57_iv_i_0[5]\, 
        edge_neg_2_sqmuxa_410_i_0, \edge_neg[4]_net_1\, 
        \edge_neg_47_iv_i_0[4]\, edge_neg_2_sqmuxa_434_i_0, 
        \edge_pos[19]_net_1\, \edge_pos_197_iv_i_0[19]\, 
        edge_pos_2_sqmuxa_402_i_0, \edge_pos[18]_net_1\, 
        \edge_pos_187_iv_i_0[18]\, N_116_0, \edge_pos[17]_net_1\, 
        \edge_pos_177_iv_i_0[17]\, edge_pos_2_sqmuxa_390_i_0, 
        \edge_pos[16]_net_1\, \edge_pos_167_iv_i_0[16]\, 
        edge_pos_2_sqmuxa_386_i_0, \edge_pos[15]_net_1\, 
        \edge_pos_157_iv_i_0[15]\, edge_pos_2_sqmuxa_404_i_0, 
        \edge_pos[14]_net_1\, \edge_pos_147_iv_i_0[14]\, 
        edge_pos_2_sqmuxa_379_i_0, \edge_pos[13]_net_1\, 
        \edge_pos_137_iv_i_0[13]\, N_216, \edge_pos[12]_net_1\, 
        N_42, \edge_pos_RNO_0[12]_net_1\, \edge_pos[11]_net_1\, 
        \edge_pos_117_iv_i_0[11]\, edge_pos_2_sqmuxa_383_i_0, 
        \edge_pos[10]_net_1\, N_44, \edge_pos_RNO_0[10]_net_1\, 
        \edge_pos[9]_net_1\, N_461_mux, N_382, 
        \edge_pos[8]_net_1\, \edge_pos_87_iv_i_0[8]\, N_36_0, 
        \edge_pos[7]_net_1\, \edge_pos_77_iv_i_0[7]\, 
        edge_pos_2_sqmuxa_387_i_0, \edge_pos[0]\, \edge_neg_7[0]\, 
        edge_pos_2_sqmuxa_i_0, \edge_neg[19]_net_1\, 
        \edge_neg_197_iv_i_0[19]\, edge_neg_2_sqmuxa_423_i_0, 
        \edge_neg[18]_net_1\, \edge_neg_187_iv_i_0[18]\, N_113_0, 
        \edge_neg[17]_net_1\, \edge_neg_177_iv_i_0[17]\, 
        edge_neg_2_sqmuxa_425_i_0, \edge_neg[16]_net_1\, 
        \edge_neg_167_iv_i_0[16]\, edge_neg_2_sqmuxa_426_i_0, 
        \edge_neg[15]_net_1\, \edge_neg_157_iv_i_0[15]\, 
        edge_neg_2_sqmuxa_427_i_0, \edge_neg[14]_net_1\, 
        \edge_neg_147_iv_i_0[14]\, edge_neg_2_sqmuxa_428_i_0, 
        \edge_neg[13]_net_1\, \edge_neg_137_iv_i_0[13]\, N_215, 
        \edge_neg[12]_net_1\, N_46, \edge_neg_RNO_0[12]_net_1\, 
        \edge_neg[11]_net_1\, \edge_neg_117_iv_i_0[11]\, 
        edge_neg_2_sqmuxa_436_i_0, \edge_neg[10]_net_1\, N_48, 
        \edge_neg_RNO_0[10]_net_1\, \edge_neg[9]_net_1\, 
        N_460_mux, N_381, \edge_neg[8]_net_1\, 
        \edge_neg_87_iv_i_0[8]\, N_37_0, \edge_neg[7]_net_1\, 
        \edge_neg_77_iv_i_0[7]\, edge_neg_2_sqmuxa_408_i_0, 
        \edge_neg[6]_net_1\, \edge_neg_67_iv_i_0[6]\, 
        edge_neg_2_sqmuxa_409_i_0, \edge_both[15]_net_1\, 
        \edge_both_157_iv_i_0[15]\, edge_both_2_sqmuxa_439_i_0, 
        \edge_both[14]_net_1\, \edge_both_147_iv_i_0[14]\, 
        edge_both_2_sqmuxa_440_i_0, \edge_both[13]_net_1\, 
        \edge_both_137_iv_i_0[13]\, N_211, \edge_both[12]_net_1\, 
        i64_mux, \edge_both_RNO_0[12]_net_1\, 
        \edge_both[11]_net_1\, \edge_both_117_iv_i_0[11]\, 
        edge_both_2_sqmuxa_452_i_0, \edge_both[10]_net_1\, 
        i15_mux, \edge_both_RNO_0[10]_net_1\, 
        \edge_both[9]_net_1\, i21_mux, \edge_both_RNO_0[9]_net_1\, 
        \edge_both[8]_net_1\, \edge_both_87_iv_i_0[8]\, N_34_0, 
        \edge_both[7]_net_1\, \edge_both_77_iv_i_0[7]\, 
        edge_both_2_sqmuxa_456_i_0, \edge_both[6]_net_1\, 
        \edge_both_67_iv_i_0[6]\, edge_both_2_sqmuxa_457_i_0, 
        \edge_both[5]_net_1\, \edge_both_57_iv_i_0[5]\, 
        edge_both_2_sqmuxa_458_i_0, \edge_both[4]_net_1\, 
        \edge_both_47_iv_i_0[4]\, edge_both_2_sqmuxa_446_i_0, 
        \edge_neg[3]\, \edge_neg_37[3]\, 
        edge_pos_2_sqmuxa_377_i_0, \edge_neg[2]\, 
        \edge_neg_27[2]\, edge_pos_2_sqmuxa_378_i_0, 
        \edge_neg[1]\, \edge_neg_17[1]\, 
        edge_pos_2_sqmuxa_399_i_0, \edge_neg[30]\, 
        \edge_neg_307[30]\, edge_pos_2_sqmuxa_391_i_0, 
        \edge_neg[29]\, \edge_neg_297[29]\, 
        edge_pos_2_sqmuxa_396_i_0, \edge_neg[28]\, 
        \edge_neg_287[28]\, edge_pos_2_sqmuxa_394_i_0, 
        \edge_neg[27]\, \edge_neg_277[27]\, 
        edge_pos_2_sqmuxa_395_i_0, \edge_pos[26]\, 
        \edge_neg_267[26]\, edge_pos_2_sqmuxa_381_i_0, 
        \edge_neg[25]\, \edge_neg_257[25]\, 
        edge_pos_2_sqmuxa_382_i_0, \edge_neg[24]\, 
        \edge_neg_247[24]\, edge_pos_2_sqmuxa_397_i_0, 
        \edge_neg[23]\, \edge_neg_237[23]\, 
        edge_pos_2_sqmuxa_398_i_0, \edge_neg[22]\, 
        \edge_neg_227[22]\, edge_pos_2_sqmuxa_392_i_0, 
        \edge_neg[21]\, \edge_neg_217[21]\, 
        edge_pos_2_sqmuxa_400_i_0, \edge_neg[20]\, 
        \edge_neg_207[20]\, edge_pos_2_sqmuxa_401_i_0, 
        \edge_both[19]_net_1\, \edge_both_197_iv_i_0[19]\, 
        edge_both_2_sqmuxa_444_i_0, \edge_both[18]_net_1\, 
        \edge_both_187_iv_i_0[18]\, N_115_0, 
        \edge_both[17]_net_1\, \edge_both_177_iv_i_0[17]\, 
        edge_both_2_sqmuxa_437_i_0, \edge_both[16]_net_1\, 
        \edge_both_167_iv_i_0[16]\, edge_both_2_sqmuxa_462_i_0, 
        \edge_neg[31]\, \edge_neg_317[31]\, edge_neg_2_sqmuxa_i_0, 
        \INTR_reg[28]_net_1\, \INTR_reg_287[28]\, 
        \INTR_reg[29]_net_1\, \INTR_reg_297[29]\, 
        \INTR_reg[30]_net_1\, \INTR_reg_307[30]\, 
        \INTR_reg[31]_net_1\, \INTR_reg_317[31]\, 
        \INTR_reg[13]_net_1\, \INTR_reg_137[13]\, 
        \INTR_reg[14]_net_1\, \INTR_reg_147[14]\, 
        \INTR_reg[15]_net_1\, \INTR_reg_157[15]\, 
        \INTR_reg[16]_net_1\, \INTR_reg_167[16]\, 
        \INTR_reg[17]_net_1\, \INTR_reg_177[17]\, 
        \INTR_reg[18]_net_1\, \INTR_reg_187[18]\, 
        \INTR_reg[19]_net_1\, \INTR_reg_197[19]\, 
        \INTR_reg[20]_net_1\, \INTR_reg_207[20]\, 
        \INTR_reg[21]_net_1\, \INTR_reg_217[21]\, 
        \INTR_reg[22]_net_1\, \INTR_reg_227[22]\, 
        \INTR_reg[23]_net_1\, \INTR_reg_237[23]\, 
        \INTR_reg[24]_net_1\, \INTR_reg_247[24]\, 
        \INTR_reg[25]_net_1\, \INTR_reg_257[25]\, 
        \INTR_reg[26]_net_1\, \INTR_reg_267[26]\, 
        \INTR_reg[27]_net_1\, \INTR_reg_277[27]\, 
        \INTR_reg[0]_net_1\, N_6172_i_0, \INTR_reg[1]_net_1\, 
        N_6167_i_0, \INTR_reg[2]_net_1\, N_6196_i_0, 
        \INTR_reg[3]_net_1\, N_6165_i_0, \INTR_reg[4]_net_1\, 
        \INTR_reg_47[4]\, \INTR_reg[5]_net_1\, N_92_i_0, 
        \INTR_reg[6]_net_1\, \INTR_reg_67[6]\, 
        \INTR_reg[7]_net_1\, N_6160_i_0, \INTR_reg[8]_net_1\, 
        \INTR_reg_87[8]\, \INTR_reg[9]_net_1\, \INTR_reg_97[9]\, 
        \INTR_reg[10]_net_1\, \INTR_reg_107[10]\, 
        \INTR_reg[11]_net_1\, \INTR_reg_117[11]\, 
        \INTR_reg[12]_net_1\, \INTR_reg_127[12]\, 
        \gpin3[6]_net_1\, \gpin2[6]_net_1\, \gpin3[7]_net_1\, 
        \gpin2[7]_net_1\, \gpin3[8]_net_1\, \gpin2[8]_net_1\, 
        \gpin3[9]_net_1\, \gpin2[9]_net_1\, \gpin3[10]_net_1\, 
        \gpin2[10]_net_1\, \gpin3[11]_net_1\, \gpin2[11]_net_1\, 
        \gpin3[12]_net_1\, \gpin2[12]_net_1\, \gpin3[13]_net_1\, 
        \gpin2[13]_net_1\, \gpin3[14]_net_1\, \gpin2[14]_net_1\, 
        \gpin3[15]_net_1\, \gpin2[15]_net_1\, \gpin3[16]_net_1\, 
        \gpin2[16]_net_1\, \gpin3[17]_net_1\, \gpin2[17]_net_1\, 
        \gpin3[18]_net_1\, \gpin2[18]_net_1\, \gpin3[19]_net_1\, 
        \gpin2[19]_net_1\, \gpin3[4]_net_1\, \gpin2[4]_net_1\, 
        \gpin3[5]_net_1\, \gpin2[5]_net_1\, \gpin1[10]_net_1\, 
        \gpin1[11]_net_1\, \gpin1[12]_net_1\, \gpin1[13]_net_1\, 
        \gpin1[14]_net_1\, \gpin1[15]_net_1\, \gpin1[16]_net_1\, 
        \gpin1[17]_net_1\, \gpin1[18]_net_1\, \gpin1[19]_net_1\, 
        \gpin1[4]_net_1\, \gpin1[5]_net_1\, \gpin1[6]_net_1\, 
        \gpin1[7]_net_1\, \gpin1[8]_net_1\, \gpin1[9]_net_1\, 
        \CONFIG_regrx[0]\, \CONFIG_regrx[1]\, \CONFIG_regrx[2]\, 
        \CONFIG_regrx[3]\, \CONFIG_regrx[4]\, \CONFIG_regrx[5]\, 
        \CONFIG_regrx[6]\, \CONFIG_regrx[7]\, CONFIG_reg_0_0_we, 
        un9_psel, m18_0, \m22_0_2\, CONFIG_rega11_2, \un30_psel\, 
        \INTR_reg_RNO_1[17]_net_1\, \INTR_reg_RNO_2[17]_net_1\, 
        N_126_0, \INTR_reg_RNO_1[14]_net_1\, 
        \INTR_reg_RNO_2[14]_net_1\, N_6250, 
        \INTR_reg_RNO_1[16]_net_1\, \INTR_reg_RNO_2[16]_net_1\, 
        N_138_0, g0_0_1_1, CONFIG_regror_9, g0_5_1, 
        CONFIG_regria_10, g0_1_2, g0_i_a3_2_0, g0_i_a3_3_0, 
        g0_i_0_1, CONFIG_regror_23_1, CONFIG_regrff_17_RNI3JFF1, 
        CONFIG_regror_10, CONFIG_rega20, g0_6_a3_0, \g0_5_0_a3_1\, 
        \g0_1_0_a3_1\, g0_6_a3_0_3, g0_6_a3_2, CONFIG_rega0, 
        CONFIG_rega4, CONFIG_regror_19, CONFIG_rega16_2, 
        CONFIG_rega9_0, g0_2_1_0, CONFIG_rega0_2, CONFIG_rega2, 
        \g0_0_1\, CONFIG_rega26_1, CONFIG_rega10, \g0_1\, 
        \g0_2_1\, CONFIG_rega21_1, CONFIG_rega1, CONFIG_rega13, 
        m23_am_1, m23_ns_1_1, m62_s_net_1, m23_ns_1, m36_am_1, 
        m36_ns_1_1, m36_ns_1, \un3_prdata_o\, m28_am_1, 
        \GPOUT_reg_RNII0ML5[6]_net_1\, m41_am_1, 
        \GPOUT_reg_RNIAKFJ5[4]_net_1\, \CONFIG_regror_29\, 
        \CONFIG_regror_28\, m52_ns_1, 
        \GPOUT_reg_RNIQ6KF5[2]_net_1\, m57_ns_1, 
        \GPOUT_reg_RNIO4KF5[1]_net_1\, CONFIG_rega18_1, 
        CONFIG_rega18, CONFIG_rega17_1, CONFIG_rega17, m62_ns_1, 
        \GPOUT_reg_RNIM2KF5[0]_net_1\, CONFIG_regria_25, 
        CONFIG_regria_23, CONFIG_regror_2, CONFIG_regror_23, 
        un15_fixed_config, m46_1, CONFIG_regror_29_1, 
        CONFIG_regror_22, CONFIG_regror_11, CONFIG_regria_31, 
        m67_0_ns_1_0, N_6195, m86_ns_1_0, N_6163, m14_ns_1, 
        N_15_0, m253_ns_1_0, N_254, m269_ns_1, N_270, m93_0_ns_1, 
        N_94_0, m239_ns_1, N_240, m161_ns_1, N_162_0, m175_ns_1, 
        N_176, m58_1_ns_1, N_59_0, m146_ns_1, N_147_0, m44_1_ns_1, 
        N_45_0, m102_ns_1_0, N_6170, \INTR_reg_RNO_1[7]_net_1\, 
        m81_ns_1, N_6158, \intr_9_u_bm[4]\, \intr_9_u_ns_1[4]\, 
        \intr_9[4]\, m20_0_ns_1, N_65, N_6243, m259_ns_1, N_257, 
        m274_ns_1, N_434_mux, \INTR_reg_227_ns_1_1[22]\, 
        \INTR_reg_227_ns_1[22]\, \INTR_reg_207_ns_1_1[20]\, 
        \INTR_reg_207_ns_1[20]\, \INTR_reg_287_ns_1_1[28]\, 
        \INTR_reg_287_ns_1[28]\, \INTR_reg_317_ns_1_1[31]\, 
        \INTR_reg_317_ns_1[31]\, \INTR_reg_277_ns_1_1[27]\, 
        \INTR_reg_277_ns_1[27]\, m99_0_ns_1, N_97_0, 
        \INTR_reg_267_ns_1_1[26]\, \INTR_reg_267_ns_1[26]\, 
        \INTR_reg_257_ns_1_1[25]\, \INTR_reg_257_ns_1[25]\, 
        \INTR_reg_307_ns_1_1[30]\, \INTR_reg_307_ns_1[30]\, 
        \INTR_reg_217_ns_1_1[21]\, \INTR_reg_217_ns_1[21]\, 
        m244_ns_1, N_433_mux, m167_ns_1, N_165_0, m50_0_ns_1, 
        N_48_0, \INTR_reg_247_ns_1_1[24]\, 
        \INTR_reg_247_ns_1[24]\, \INTR_reg_237_ns_1_1[23]\, 
        \INTR_reg_237_ns_1[23]\, m181_ns_1, N_179, m64_1_ns_1, 
        N_62_0, m152_ns_1, N_150_0, \INTR_reg_297_ns_1_1[29]\, 
        \INTR_reg_297_ns_1[29]\, m309_ns_1, m332_ns_1, m337_ns_1, 
        m342_ns_1, m318_ns_1, \N_6186\, m323_ns_1, m352_ns_1, 
        m357_ns_1, m327_ns_1, un249_fixed_config, 
        un977_fixed_config, un957_fixed_config, 
        un229_fixed_config, un1107_fixed_config, 
        un659_fixed_config, un883_fixed_config, 
        un379_fixed_config, un939_fixed_config, 
        un921_fixed_config, un901_fixed_config, 
        un995_fixed_config, un267_fixed_config, un1_psel_280_2, 
        un789_fixed_config, un809_fixed_config, 
        un827_fixed_config, CONFIG_rega12_1, CONFIG_rega23_2, 
        \CONFIG_rega23_1\, CONFIG_rega25_2, CONFIG_rega26_2, 
        CONFIG_rega30_2, CONFIG_rega30_1, N_6193, N_5144, 
        CONFIG_regria_5_0, CONFIG_regria_24_0, CONFIG_regria_8_0, 
        CONFIG_rega8_0, CONFIG_rega0_0, CONFIG_rega3_0, 
        CONFIG_rega28_0, CONFIG_rega22_0, CONFIG_rega30_0, 
        CONFIG_rega24_0, CONFIG_rega16_0, CONFIG_rega21_0, 
        CONFIG_rega29_0, CONFIG_rega25_0, CONFIG_rega5_0, N_6155, 
        N_70, N_6152, N_22_0, N_25_0, N_6244, N_75_0, N_101_0, 
        N_104_0, N_186, N_195, N_201, N_279, N_285, N_296, N_198, 
        N_192, N_189, N_183, N_107_0, N_377, N_374, N_288, N_72_0, 
        N_66_0, N_69_0, N_6191, N_6192, N_6190, N_292, N_282, 
        N_276, N_88, CONFIG_rega7, CONFIG_rega6, CONFIG_rega26, 
        CONFIG_regria_30, CONFIG_regria_29, CONFIG_regria_28, 
        CONFIG_regria_27, CONFIG_regria_22, CONFIG_regria_21, 
        CONFIG_regria_16, CONFIG_regria_15, CONFIG_regria_12, 
        CONFIG_regria_3, N_6174, N_6177, CONFIG_regror_0, 
        CONFIG_regria_26, CONFIG_regria_19, CONFIG_regria_11, 
        \intr_7[3]\, \intr_3[1]\, CONFIG_regror_18, 
        CONFIG_regror_17, CONFIG_regror_16, un11_psel_1_0, N_90
         : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc28, nc14, nc5, nc21, nc15, nc3, nc10, nc7, 
        nc17, nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11
         : std_logic;

begin 

    GPOUT_reg_31 <= \GPOUT_reg_31\;
    un30_psel <= \un30_psel\;
    m62_s <= m62_s_net_1;
    un3_prdata_o <= \un3_prdata_o\;
    CONFIG_regror_29 <= \CONFIG_regror_29\;
    CONFIG_regror_28 <= \CONFIG_regror_28\;
    N_6186 <= \N_6186\;
    CONFIG_rega23_1 <= \CONFIG_rega23_1\;

    \CONFIG_reg_5_RNILD2U2[1]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => \INTR_reg[5]_net_1\, B => 
        \CONFIG_reg_5[1]_net_1\, C => \un3_prdata_o\, D => 
        \gpin3[5]_net_1\, Y => m36_am_1);
    
    edge_both_2_sqmuxa_437_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_17[3]_net_1\, D => un995_fixed_config, Y => 
        edge_both_2_sqmuxa_437_i_0);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIMRH78\ : 
        CFG4
      generic map(INIT => x"2075")

      port map(A => m62_s_net_1, B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => \CONFIG_regrx[0]\, D
         => \GPOUT_reg_RNIM2KF5[0]_net_1\, Y => m62_ns_1);
    
    \edge_pos[7]\ : SLE
      port map(D => \edge_pos_77_iv_i_0[7]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_387_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[7]_net_1\);
    
    \CONFIG_reg_1[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un41_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_1[5]_net_1\);
    
    \GPOUT_reg[15]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(15), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[15]_net_1\);
    
    \GEN_BITS.21.APB_32.INTR_reg_217_ns_1_1[21]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_21[5]_net_1\, B => \edge_neg[21]\, 
        C => \CONFIG_reg_21[7]_net_1\, D => 
        \CONFIG_reg_21[6]_net_1\, Y => \INTR_reg_217_ns_1_1[21]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_13\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un387_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_13);
    
    edge_pos_2_sqmuxa_388_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[6]_net_1\, B => N_65, C => 
        \gpin3[6]_net_1\, D => \CONFIG_reg_6[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_388_i_0);
    
    \INTR_reg_RNO_3[13]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_13[6]_net_1\, B => 
        \edge_pos[13]_net_1\, C => \gpin3[13]_net_1\, D => 
        \CONFIG_reg_13[7]_net_1\, Y => m161_ns_1);
    
    \CONFIG_reg_18[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un532_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_18[7]_net_1\);
    
    \edge_pos[11]\ : SLE
      port map(D => \edge_pos_117_iv_i_0[11]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_383_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[11]_net_1\);
    
    \GEN_BITS.17.APB_32.un995_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[17]_net_1\, B => \gpin3[17]_net_1\, Y
         => un995_fixed_config);
    
    \GPOUT_reg[25]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(25), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_25);
    
    \gpin1[17]\ : SLE
      port map(D => GPIO_IN_c(17), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[17]_net_1\);
    
    \CONFIG_reg_27[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un793_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_27[6]_net_1\);
    
    \edge_neg[19]\ : SLE
      port map(D => \edge_neg_197_iv_i_0[19]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_423_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[19]_net_1\);
    
    \GEN_BITS.20.APB_32.INTR_reg_207_ns[20]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(20), B => N_65, 
        C => \INTR_reg[20]_net_1\, D => \INTR_reg_207_ns_1[20]\, 
        Y => \INTR_reg_207[20]\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_5\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega30_2, B => CONFIG_rega29_0, C => 
        un9_psel, D => m18_0, Y => un851_psel);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_22\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega0, Y
         => un11_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_31_RNI926M6\ : CFG3
      generic map(INIT => x"01")

      port map(A => CONFIG_regror_10, B => CONFIG_regria_31, C
         => CONFIG_regror_9, Y => CONFIG_regror_29_1);
    
    \CONFIG_reg_18[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un532_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_18[6]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_23_RNI2N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega23_2, B => \CONFIG_rega23_1\, C
         => CONFIG_regro_23, D => CoreAPB3_0_APBmslave0_PADDR(5), 
        Y => CONFIG_regria_23);
    
    \CONFIG_reg_24[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un706_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_24[5]_net_1\);
    
    \edge_both_RNO[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[1]\, B => \CONFIG_reg_1[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(1), Y => 
        \edge_neg_17[1]\);
    
    \edge_pos_RNO[9]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[9]_net_1\, B => N_377, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        N_461_mux);
    
    \GEN_BITS.17.APB_32.un957_fixed_config\ : CFG2
      generic map(INIT => x"2")

      port map(A => \gpin2[17]_net_1\, B => \gpin3[17]_net_1\, Y
         => un957_fixed_config);
    
    \gpin2[12]\ : SLE
      port map(D => \gpin1[12]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[12]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega0_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega0_0);
    
    \GPOUT_reg_RNIO4KF5[1]\ : CFG4
      generic map(INIT => x"23EF")

      port map(A => \un3_prdata_o\, B => \un30_psel\, C => 
        \INTR_reg[1]_net_1\, D => \GPOUT_reg[1]_net_1\, Y => 
        \GPOUT_reg_RNIO4KF5[1]_net_1\);
    
    \gpin1[5]\ : SLE
      port map(D => GPIO_IN_c(5), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[5]_net_1\);
    
    \edge_pos[16]\ : SLE
      port map(D => \edge_pos_167_iv_i_0[16]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_386_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[16]_net_1\);
    
    \GEN_BITS.31.APB_32.INTR_reg_317_ns_1_1[31]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_31[5]_net_1\, B => \edge_neg[31]\, 
        C => \CONFIG_reg_31[7]_net_1\, D => 
        \CONFIG_reg_31[6]_net_1\, Y => \INTR_reg_317_ns_1_1[31]\);
    
    \CONFIG_reg_28[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un822_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_28[5]_net_1\);
    
    \INTR_reg_RNISL6H2[28]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[28]_net_1\, Y => N_440);
    
    \CONFIG_reg_27[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un793_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_27[3]_net_1\);
    
    \GEN_BITS.27.APB_32.INTR_reg_277_ns[27]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(27), B => N_65, 
        C => \INTR_reg[27]_net_1\, D => \INTR_reg_277_ns_1[27]\, 
        Y => \INTR_reg_277[27]\);
    
    \GPOUT_reg_RNIEIQ752[7]\ : CFG4
      generic map(INIT => x"3373")

      port map(A => \CONFIG_regror_29\, B => m23_ns_1, C => 
        m62_s_net_1, D => \CONFIG_regror_28\, Y => N_24_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_2_RNI51BA1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => CONFIG_regro_2, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => g0_6_a3_0_3);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_14\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un416_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_14);
    
    \edge_both_RNO_0[30]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_30[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_391_i_0);
    
    \CONFIG_reg_25[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un735_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_25[5]_net_1\);
    
    \CONFIG_reg_0[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un11_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_0[6]_net_1\);
    
    \CONFIG_reg_21[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un619_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_21[3]_net_1\);
    
    \GEN_BITS.15.APB_32.edge_both_157_iv_i[15]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[15]_net_1\, B => 
        \CONFIG_reg_15[3]_net_1\, C => un883_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(15), Y => 
        \edge_both_157_iv_i_0[15]\);
    
    \GPOUT_reg_RNIM2KF5[0]\ : CFG4
      generic map(INIT => x"2E3F")

      port map(A => \un3_prdata_o\, B => \un30_psel\, C => 
        \GPOUT_reg[0]_net_1\, D => \INTR_reg[0]_net_1\, Y => 
        \GPOUT_reg_RNIM2KF5[0]_net_1\);
    
    \edge_neg_RNO_1[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[10]_net_1\, B => 
        \CONFIG_reg_10[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(10), Y => N_276);
    
    \INTR_reg_RNO_2[9]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \edge_both[9]_net_1\, B => 
        \CONFIG_reg_9[5]_net_1\, C => \CONFIG_reg_9[6]_net_1\, D
         => \CONFIG_reg_9[3]_net_1\, Y => N_433_mux);
    
    \INTR_reg_RNO_0[6]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_6[7]_net_1\, B => 
        \CONFIG_reg_6[5]_net_1\, C => N_45_0, D => N_48_0, Y => 
        m50_0_ns_1);
    
    \edge_both_RNO[18]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[18]_net_1\, B => N_65, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        N_115_0);
    
    \INTR_reg_RNO_0[18]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_18[7]_net_1\, B => 
        \CONFIG_reg_18[5]_net_1\, C => N_94_0, D => N_97_0, Y => 
        m99_0_ns_1);
    
    \gpin1[7]\ : SLE
      port map(D => GPIO_IN_c(7), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[7]_net_1\);
    
    \CONFIG_reg_6_RNIOI5V2[1]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => \INTR_reg[6]_net_1\, B => 
        \CONFIG_reg_6[1]_net_1\, C => \un3_prdata_o\, D => 
        \gpin3[6]_net_1\, Y => m28_am_1);
    
    \INTR_reg[30]\ : SLE
      port map(D => \INTR_reg_307[30]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[30]_net_1\);
    
    \gpin1[15]\ : SLE
      port map(D => GPIO_IN_c(15), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[15]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega30_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => CONFIG_rega30_0);
    
    \GEN_BITS.8.APB_32.edge_both_87_iv_i_RNO[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[8]_net_1\, B => 
        \CONFIG_reg_8[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(8), Y => N_6244);
    
    \GEN_BITS.13.APB_32.edge_pos_137_iv_i[13]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[13]_net_1\, B => N_195, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        \edge_pos_137_iv_i_0[13]\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_16\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega6, Y
         => un185_psel);
    
    \INTR_reg_RNO[10]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[10]_net_1\, B => m259_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(10), D => N_65, Y => 
        \INTR_reg_107[10]\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNI8IP45_0\ : 
        CFG4
      generic map(INIT => x"0C55")

      port map(A => \un30_psel\, B => \CONFIG_regrx[7]\, C => 
        CoreAPB3_0_APBmslave0_PADDR(7), D => m62_s_net_1, Y => 
        m23_ns_1_1);
    
    \CONFIG_reg_30[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un880_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_30[3]_net_1\);
    
    \CONFIG_reg_0[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un11_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_0[3]_net_1\);
    
    \gpin2[4]\ : SLE
      port map(D => \gpin1[4]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[4]_net_1\);
    
    \CONFIG_reg_6[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un185_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_6[1]_net_1\);
    
    \edge_pos_RNO[12]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[12]_net_1\, B => N_285, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        N_42);
    
    \edge_both[5]\ : SLE
      port map(D => \edge_both_57_iv_i_0[5]\, CLK => FAB_CCC_GL0, 
        EN => edge_both_2_sqmuxa_458_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[5]_net_1\);
    
    \GEN_BITS.30.APB_32.INTR_reg_307_ns[30]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(30), B => N_65, 
        C => \INTR_reg[30]_net_1\, D => \INTR_reg_307_ns_1[30]\, 
        Y => \INTR_reg_307[30]\);
    
    \INTR_reg_RNO_2[13]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[13]_net_1\, B => 
        \CONFIG_reg_13[3]_net_1\, C => \edge_neg[13]_net_1\, D
         => \CONFIG_reg_13[6]_net_1\, Y => N_165_0);
    
    \INTR_reg_RNO_0[12]\ : CFG3
      generic map(INIT => x"2E")

      port map(A => N_270, B => \CONFIG_reg_12[7]_net_1\, C => 
        N_434_mux, Y => m274_ns_1);
    
    \INTR_reg[29]\ : SLE
      port map(D => \INTR_reg_297[29]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[29]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIDNDGT1\ : 
        CFG4
      generic map(INIT => x"54AA")

      port map(A => un15_fixed_config, B => \CONFIG_regror_28\, C
         => \CONFIG_regror_29\, D => m46_1, Y => N_47);
    
    \CONFIG_reg_26[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un764_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_26[5]_net_1\);
    
    \CONFIG_reg_25[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un735_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_25[7]_net_1\);
    
    \GPOUT_reg_RNI36165[9]\ : CFG4
      generic map(INIT => x"15BF")

      port map(A => \N_6186\, B => \un30_psel\, C => 
        \GPOUT_reg[9]_net_1\, D => \INTR_reg[9]_net_1\, Y => 
        m352_ns_1);
    
    \INTR_reg_RNO_2[6]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[6]_net_1\, B => 
        \CONFIG_reg_6[3]_net_1\, C => \edge_neg[6]_net_1\, D => 
        \CONFIG_reg_6[6]_net_1\, Y => N_48_0);
    
    \INTR_reg[18]\ : SLE
      port map(D => \INTR_reg_187[18]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[18]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_17\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega7, Y
         => un214_psel);
    
    \GEN_BITS.21.APB_32.INTR_reg_217_ns_1[21]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_217_ns_1_1[21]\, B => 
        \CONFIG_reg_21[3]_net_1\, Y => \INTR_reg_217_ns_1[21]\);
    
    \edge_neg[12]\ : SLE
      port map(D => N_46, CLK => FAB_CCC_GL0, EN => 
        \edge_neg_RNO_0[12]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[12]_net_1\);
    
    \CONFIG_reg_1[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un41_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_1[7]_net_1\);
    
    \edge_both_RNO[24]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[24]\, B => \CONFIG_reg_24[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(24), Y => 
        \edge_neg_247[24]\);
    
    \GEN_BITS.4.REG_INT.intr_9_u_ns[4]\ : CFG4
      generic map(INIT => x"A820")

      port map(A => \CONFIG_reg_4[3]_net_1\, B => 
        \CONFIG_reg_4[7]_net_1\, C => \intr_9_u_bm[4]\, D => 
        \intr_9_u_ns_1[4]\, Y => \intr_9[4]\);
    
    \GEN_BITS.15.APB_32.un883_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[15]_net_1\, B => \gpin3[15]_net_1\, Y
         => un883_fixed_config);
    
    \edge_both_RNO[0]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[0]\, B => \CONFIG_reg_0[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(0), Y => 
        \edge_neg_7[0]\);
    
    \gpin3[10]\ : SLE
      port map(D => \gpin2[10]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[10]_net_1\);
    
    \gpin1[6]\ : SLE
      port map(D => GPIO_IN_c(6), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[6]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNI8IP45\ : 
        CFG4
      generic map(INIT => x"0C55")

      port map(A => \un30_psel\, B => \CONFIG_regrx[5]\, C => 
        CoreAPB3_0_APBmslave0_PADDR(7), D => m62_s_net_1, Y => 
        m36_ns_1_1);
    
    \CONFIG_reg_29[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un851_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_29[7]_net_1\);
    
    \edge_both_RNO_0[1]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_1[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_399_i_0);
    
    \edge_both[30]\ : SLE
      port map(D => \edge_neg_307[30]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_391_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[30]\);
    
    \CONFIG_reg_26[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un764_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_26[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega22_0\ : CFG3
      generic map(INIT => x"20")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega22_0);
    
    \CONFIG_reg_22[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un648_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_22[3]_net_1\);
    
    \CONFIG_reg_20[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un590_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_20[6]_net_1\);
    
    edge_both_2_sqmuxa_462_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_16[3]_net_1\, D => un939_fixed_config, Y => 
        edge_both_2_sqmuxa_462_i_0);
    
    \INTR_reg_RNO[17]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[17]_net_1\, B => N_126_0, C => 
        CoreAPB3_0_APBmslave0_PWDATA(17), D => N_65, Y => 
        \INTR_reg_177[17]\);
    
    \INTR_reg_RNO_2[16]\ : CFG4
      generic map(INIT => x"5066")

      port map(A => \CONFIG_reg_16[5]_net_1\, B => 
        \gpin3[16]_net_1\, C => \edge_both[16]_net_1\, D => 
        \CONFIG_reg_16[7]_net_1\, Y => \INTR_reg_RNO_2[16]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_1_RNIM9MB2\ : CFG4
      generic map(INIT => x"0002")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => g0_0_1_1, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_regror_9);
    
    \INTR_reg_RNIMF6H2[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[22]_net_1\, Y => INTR_reg_m_0);
    
    \gpin3[8]\ : SLE
      port map(D => \gpin2[8]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[8]_net_1\);
    
    \INTR_reg_RNO_1[5]\ : CFG4
      generic map(INIT => x"35FF")

      port map(A => \edge_pos[5]_net_1\, B => \edge_neg[5]_net_1\, 
        C => \CONFIG_reg_5[5]_net_1\, D => 
        \CONFIG_reg_5[3]_net_1\, Y => N_88);
    
    \INTR_reg_RNILE6H2[21]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[21]_net_1\, Y => N_437);
    
    \GEN_BITS.8.APB_32.edge_pos_87_iv_i_RNO[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[8]_net_1\, B => 
        \CONFIG_reg_8[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(8), Y => N_25_0);
    
    \CONFIG_reg_20[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un590_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_20[7]_net_1\);
    
    \GEN_BITS.5.APB_32.edge_neg_57_iv_i_RNO[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[5]_net_1\, B => 
        \CONFIG_reg_5[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(5), Y => N_6155);
    
    \GPOUT_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[2]_net_1\);
    
    \gpin3[18]\ : SLE
      port map(D => \gpin2[18]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[18]_net_1\);
    
    \GEN_BITS.4.APB_32.INTR_reg_47[4]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => N_65, C
         => \INTR_reg[4]_net_1\, D => \intr_9[4]\, Y => 
        \INTR_reg_47[4]\);
    
    g0_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => \g0_0_1\, Y => 
        CONFIG_rega10);
    
    \CONFIG_reg_8_RNIKP78[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \gpin3[8]_net_1\, B => 
        \CONFIG_reg_8[1]_net_1\, Y => N_426_mux);
    
    \CONFIG_reg_27[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un793_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_27[7]_net_1\);
    
    edge_neg_2_sqmuxa_410_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[5]_net_1\, B => N_65, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_410_i_0);
    
    \edge_neg[18]\ : SLE
      port map(D => \edge_neg_187_iv_i_0[18]\, CLK => FAB_CCC_GL0, 
        EN => N_113_0, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_neg[18]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_14_RNI88TU2\ : CFG4
      generic map(INIT => x"EC00")

      port map(A => CONFIG_regro_14, B => CONFIG_regria_8_0, C
         => CONFIG_rega30_1, D => CONFIG_rega8_0, Y => 
        CONFIG_regror_0);
    
    \GEN_BITS.4.APB_32.edge_neg_47_iv_i[4]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_neg[4]_net_1\, B => 
        \CONFIG_reg_4[3]_net_1\, C => un249_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(4), Y => 
        \edge_neg_47_iv_i_0[4]\);
    
    g0_6 : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega26_1);
    
    \edge_both[14]\ : SLE
      port map(D => \edge_both_147_iv_i_0[14]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_440_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[14]_net_1\);
    
    \INTR_reg[14]\ : SLE
      port map(D => \INTR_reg_147[14]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[14]_net_1\);
    
    \GPOUT_reg_RNIVIG25[16]\ : CFG4
      generic map(INIT => x"15BF")

      port map(A => \N_6186\, B => \un30_psel\, C => 
        \GPOUT_reg[16]_net_1\, D => \INTR_reg[16]_net_1\, Y => 
        m327_ns_1);
    
    \CONFIG_reg_22[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un648_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_22[5]_net_1\);
    
    \gpin2[11]\ : SLE
      port map(D => \gpin1[11]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[11]_net_1\);
    
    \GEN_BITS.13.APB_32.edge_pos_137_iv_i_RNO[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[13]_net_1\, B => 
        \CONFIG_reg_13[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(13), Y => N_195);
    
    \GEN_BITS.15.APB_32.edge_neg_157_iv_i_RNO[15]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[15]_net_1\, B => 
        \CONFIG_reg_15[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(15), Y => N_189);
    
    \CONFIG_reg_8[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un242_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_8[3]_net_1\);
    
    \GPOUT_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[0]_net_1\);
    
    \GEN_BITS.23.APB_32.INTR_reg_237_ns_1[23]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_237_ns_1_1[23]\, B => 
        \CONFIG_reg_23[3]_net_1\, Y => \INTR_reg_237_ns_1[23]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega12_1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega12_1);
    
    \edge_pos[12]\ : SLE
      port map(D => N_42, CLK => FAB_CCC_GL0, EN => 
        \edge_pos_RNO_0[12]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[12]_net_1\);
    
    \edge_both_RNO[8]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[8]_net_1\, B => N_65, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        N_34_0);
    
    \edge_both[23]\ : SLE
      port map(D => \edge_neg_237[23]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_398_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[23]\);
    
    \CONFIG_reg_27[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un793_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_27[5]_net_1\);
    
    \gpin1[19]\ : SLE
      port map(D => GPIO_IN_c(19), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[19]_net_1\);
    
    \CONFIG_reg_25[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un735_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_25[6]_net_1\);
    
    \CONFIG_reg_16[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un474_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_16[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \INTR_reg_RNO[12]\ : CFG4
      generic map(INIT => x"330A")

      port map(A => \INTR_reg[12]_net_1\, B => m274_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(12), D => N_65, Y => 
        \INTR_reg_127[12]\);
    
    \INTR_reg[22]\ : SLE
      port map(D => \INTR_reg_227[22]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[22]_net_1\);
    
    \INTR_reg_RNO_1[18]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_18[3]_net_1\, B => m93_0_ns_1, C
         => \edge_both[18]_net_1\, D => \CONFIG_reg_18[7]_net_1\, 
        Y => N_94_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_30\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un880_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_30);
    
    \edge_neg[6]\ : SLE
      port map(D => \edge_neg_67_iv_i_0[6]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_409_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[6]_net_1\);
    
    \CONFIG_reg_6[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un185_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_6[6]_net_1\);
    
    \INTR_reg_RNO[14]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[14]_net_1\, B => N_6250, C => 
        CoreAPB3_0_APBmslave0_PWDATA(14), D => N_65, Y => 
        \INTR_reg_147[14]\);
    
    \gpin3[4]\ : SLE
      port map(D => \gpin2[4]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[4]_net_1\);
    
    \GEN_BITS.16.APB_32.edge_neg_167_iv_i[16]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_neg[16]_net_1\, B => 
        \CONFIG_reg_16[3]_net_1\, C => un921_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(16), Y => 
        \edge_neg_167_iv_i_0[16]\);
    
    \CONFIG_reg_14[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un416_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_14[3]_net_1\);
    
    \GEN_BITS.16.APB_32.un921_fixed_config\ : CFG2
      generic map(INIT => x"4")

      port map(A => \gpin2[16]_net_1\, B => \gpin3[16]_net_1\, Y
         => un921_fixed_config);
    
    \INTR_reg_RNO[19]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[19]_net_1\, B => m64_1_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(19), D => N_65, Y => 
        \INTR_reg_197[19]\);
    
    \CONFIG_reg_7[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un214_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_7[7]_net_1\);
    
    \CONFIG_reg_22[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un648_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_22[7]_net_1\);
    
    \edge_pos_RNO_1[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[10]_net_1\, B => 
        \CONFIG_reg_10[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(10), Y => N_282);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega25_2, B => CONFIG_rega21_0, C => 
        un9_psel, D => m18_0, Y => un619_psel);
    
    \INTR_reg_RNIQJ6H2[26]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[26]_net_1\, Y => INTR_reg_m_4);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_0_RNIAKDL3\ : CFG4
      generic map(INIT => x"1110")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => g0_6_a3_0_3, D => 
        g0_6_a3_2, Y => CONFIG_regror_19);
    
    \CONFIG_reg_4[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un127_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_4[1]_net_1\);
    
    \INTR_reg_RNO[3]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => N_65, C
         => \INTR_reg[3]_net_1\, D => \intr_7[3]\, Y => 
        N_6165_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_23\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un677_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_23);
    
    \CONFIG_reg_13[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un387_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_13[3]_net_1\);
    
    \CONFIG_reg_9[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un271_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_9[6]_net_1\);
    
    \INTR_reg[26]\ : SLE
      port map(D => \INTR_reg_267[26]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[26]_net_1\);
    
    \GPOUT_reg_RNIUOIRA[7]\ : CFG4
      generic map(INIT => x"CC74")

      port map(A => m23_am_1, B => m23_ns_1_1, C => 
        \GPOUT_reg[7]_net_1\, D => m62_s_net_1, Y => m23_ns_1);
    
    \gpin2[8]\ : SLE
      port map(D => \gpin1[8]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[8]_net_1\);
    
    \CONFIG_reg_2[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un69_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_2[5]_net_1\);
    
    \INTR_reg_RNO_1[12]\ : CFG4
      generic map(INIT => x"D7DD")

      port map(A => \CONFIG_reg_12[3]_net_1\, B => m269_ns_1, C
         => \CONFIG_reg_12[6]_net_1\, D => \gpin3[12]_net_1\, Y
         => N_270);
    
    \GPOUT_reg[16]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(16), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[16]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_12_RNIE3HQ5\ : CFG3
      generic map(INIT => x"FE")

      port map(A => CONFIG_regria_19, B => CONFIG_regria_12, C
         => CONFIG_regria_28, Y => CONFIG_regror_17);
    
    \edge_pos[9]\ : SLE
      port map(D => N_461_mux, CLK => FAB_CCC_GL0, EN => N_382, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \edge_pos[9]_net_1\);
    
    \CONFIG_reg_14[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un416_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_14[1]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega23_1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \CONFIG_rega23_1\);
    
    \GEN_BITS.13.APB_32.edge_neg_137_iv_i[13]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[13]_net_1\, B => N_186, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        \edge_neg_137_iv_i_0[13]\);
    
    \INTR_reg_RNO_0[13]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_13[7]_net_1\, B => 
        \CONFIG_reg_13[5]_net_1\, C => N_162_0, D => N_165_0, Y
         => m167_ns_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_15\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CONFIG_rega12_1, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un445_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_18\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un532_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_18);
    
    \INTR_reg_RNO_1[6]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_6[3]_net_1\, B => m44_1_ns_1, C
         => \edge_both[6]_net_1\, D => \CONFIG_reg_6[7]_net_1\, Y
         => N_45_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega26\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => CONFIG_rega26_1, D
         => CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega26);
    
    \INTR_reg_RNO_3[10]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \CONFIG_reg_10[7]_net_1\, B => 
        \edge_both[10]_net_1\, C => \CONFIG_reg_10[5]_net_1\, Y
         => m253_ns_1_0);
    
    \edge_pos_RNO_1[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[12]_net_1\, B => 
        \CONFIG_reg_12[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(12), Y => N_285);
    
    \GPOUT_reg[26]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(26), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_26);
    
    \INTR_reg_RNO_3[5]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \CONFIG_reg_5[7]_net_1\, B => 
        \edge_both[5]_net_1\, C => \CONFIG_reg_5[5]_net_1\, Y => 
        m86_ns_1_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_15_RNI3M5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega12_1, B => \CONFIG_rega23_1\, C
         => CONFIG_regro_15, D => CoreAPB3_0_APBmslave0_PADDR(6), 
        Y => CONFIG_regria_15);
    
    \CONFIG_reg_21[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un619_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_21[5]_net_1\);
    
    \gpin2[13]\ : SLE
      port map(D => \gpin1[13]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[13]_net_1\);
    
    \GEN_BITS.6.APB_32.un379_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[6]_net_1\, B => \gpin3[6]_net_1\, Y
         => un379_fixed_config);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_24\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un706_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_24);
    
    \CONFIG_reg_21[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un619_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_21[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega17_1\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega17_1);
    
    \CONFIG_reg_19_RNIA6G78[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_19[1]_net_1\, B => 
        \gpin3[19]_net_1\, C => \un3_prdata_o\, D => m342_ns_1, Y
         => N_343);
    
    \edge_both_RNO_0[22]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_22[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_392_i_0);
    
    \INTR_reg_RNO_0[16]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \CONFIG_reg_16[6]_net_1\, B => 
        \CONFIG_reg_16[3]_net_1\, C => \INTR_reg_RNO_1[16]_net_1\, 
        D => \INTR_reg_RNO_2[16]_net_1\, Y => N_138_0);
    
    \INTR_reg_RNO_2[5]\ : CFG4
      generic map(INIT => x"8882")

      port map(A => \CONFIG_reg_5[3]_net_1\, B => m86_ns_1_0, C
         => \CONFIG_reg_5[7]_net_1\, D => \gpin3[5]_net_1\, Y => 
        N_6163);
    
    \GEN_BITS.16.APB_32.edge_pos_167_iv_i[16]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_pos[16]_net_1\, B => 
        \CONFIG_reg_16[3]_net_1\, C => un901_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(16), Y => 
        \edge_pos_167_iv_i_0[16]\);
    
    \edge_both[2]\ : SLE
      port map(D => \edge_neg_27[2]\, CLK => FAB_CCC_GL0, EN => 
        edge_pos_2_sqmuxa_378_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[2]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega26_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => CONFIG_rega26_2);
    
    \GPOUT_reg_RNIJ6G25[10]\ : CFG4
      generic map(INIT => x"15BF")

      port map(A => \N_6186\, B => \un30_psel\, C => 
        \GPOUT_reg[10]_net_1\, D => \INTR_reg[10]_net_1\, Y => 
        m357_ns_1);
    
    \INTR_reg_RNO[18]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[18]_net_1\, B => m99_0_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(18), D => N_65, Y => 
        \INTR_reg_187[18]\);
    
    \edge_pos[6]\ : SLE
      port map(D => \edge_pos_67_iv_i_0[6]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_388_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[6]_net_1\);
    
    \INTR_reg_RNO_0[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_6174, B => \CONFIG_reg_3[3]_net_1\, Y => 
        \intr_7[3]\);
    
    \edge_neg_RNO_1[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[12]_net_1\, B => 
        \CONFIG_reg_12[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(12), Y => N_279);
    
    \GEN_BITS.18.APB_32.edge_neg_187_iv_i_RNO[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[18]_net_1\, B => 
        \CONFIG_reg_18[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(18), Y => N_101_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_22_RNI1N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega30_1, B => CONFIG_rega26_2, C => 
        CONFIG_regro_22, D => CoreAPB3_0_APBmslave0_PADDR(5), Y
         => CONFIG_regria_22);
    
    \INTR_reg[17]\ : SLE
      port map(D => \INTR_reg_177[17]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[17]_net_1\);
    
    \INTR_reg_RNO_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => m102_ns_1_0, B => \CONFIG_reg_0[3]_net_1\, Y
         => N_6170);
    
    \INTR_reg[15]\ : SLE
      port map(D => \INTR_reg_157[15]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[15]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_17\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un503_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_17);
    
    \INTR_reg_RNIMG7H2[31]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[31]_net_1\, Y => INTR_reg_m_9);
    
    \edge_neg[4]\ : SLE
      port map(D => \edge_neg_47_iv_i_0[4]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_434_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[4]_net_1\);
    
    \CONFIG_reg_23[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un677_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_23[6]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_21_RNI9TMO7\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => CONFIG_regria_29, B => CONFIG_regria_22, C
         => CONFIG_regria_21, D => CONFIG_regria_30, Y => 
        CONFIG_regror_16);
    
    \GPOUT_reg_RNIQ6KF5[2]\ : CFG4
      generic map(INIT => x"23EF")

      port map(A => \un3_prdata_o\, B => \un30_psel\, C => 
        \INTR_reg[2]_net_1\, D => \GPOUT_reg[2]_net_1\, Y => 
        \GPOUT_reg_RNIQ6KF5[2]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNITT543\ : 
        CFG4
      generic map(INIT => x"0A4E")

      port map(A => un15_fixed_config, B => \CONFIG_regrx[3]\, C
         => \INTR_reg[3]_net_1\, D => 
        CoreAPB3_0_APBmslave0_PADDR(7), Y => m46_1);
    
    \edge_both_RNO_0[31]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_31[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_neg_2_sqmuxa_i_0);
    
    \GEN_BITS.20.APB_32.INTR_reg_207_ns_1[20]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_207_ns_1_1[20]\, B => 
        \CONFIG_reg_20[3]_net_1\, Y => \INTR_reg_207_ns_1[20]\);
    
    \GEN_BITS.7.APB_32.edge_pos_77_iv_i[7]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[7]_net_1\, B => N_6191, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        \edge_pos_77_iv_i_0[7]\);
    
    \edge_both_RNO[9]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[9]_net_1\, B => N_288, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        i21_mux);
    
    \CONFIG_reg_16[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un474_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_16[3]_net_1\);
    
    \INTR_reg_RNO[15]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[15]_net_1\, B => m181_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(15), D => N_65, Y => 
        \INTR_reg_157[15]\);
    
    \CONFIG_reg_19[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un561_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_19[3]_net_1\);
    
    \CONFIG_reg_13[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un387_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_13[5]_net_1\);
    
    \GEN_BITS.4.REG_INT.intr_9_1[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \edge_pos[4]_net_1\, B => \edge_neg[4]_net_1\, 
        C => \CONFIG_reg_4[5]_net_1\, Y => N_5144);
    
    \INTR_reg_RNO_2[10]\ : CFG4
      generic map(INIT => x"35FF")

      port map(A => \edge_pos[10]_net_1\, B => 
        \edge_neg[10]_net_1\, C => \CONFIG_reg_10[5]_net_1\, D
         => \CONFIG_reg_10[3]_net_1\, Y => N_257);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_7\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega30_2, B => CONFIG_rega30_0, C => 
        un9_psel, D => m18_0, Y => un880_psel);
    
    \INTR_reg_RNO[11]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[11]_net_1\, B => m152_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(11), D => N_65, Y => 
        \INTR_reg_117[11]\);
    
    \CONFIG_reg_31[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un909_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_31[3]_net_1\);
    
    \GEN_BITS.5.APB_32.edge_pos_57_iv_i_RNO[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[5]_net_1\, B => 
        \CONFIG_reg_5[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(5), Y => N_70);
    
    edge_neg_2_sqmuxa_436_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[11]_net_1\, B => N_65, C => 
        \gpin3[11]_net_1\, D => \CONFIG_reg_11[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_436_i_0);
    
    \INTR_reg_RNO_2[7]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \edge_both[7]_net_1\, B => 
        \CONFIG_reg_7[6]_net_1\, C => \CONFIG_reg_7[5]_net_1\, Y
         => m81_ns_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_8_RNI6IN01\ : CFG3
      generic map(INIT => x"02")

      port map(A => CONFIG_regro_8, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_regria_8_0);
    
    edge_both_2_sqmuxa_446_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_4[3]_net_1\, D => un267_fixed_config, Y => 
        edge_both_2_sqmuxa_446_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_20_RNILOUA1\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => CONFIG_regro_20, D
         => CoreAPB3_0_APBmslave0_PADDR(4), Y => g0_i_0_1);
    
    \CONFIG_reg_10[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un300_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_10[5]_net_1\);
    
    \GPOUT_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[4]_net_1\);
    
    \INTR_reg_RNO_3[8]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_8[6]_net_1\, B => 
        \edge_pos[8]_net_1\, C => \gpin3[8]_net_1\, D => 
        \CONFIG_reg_8[7]_net_1\, Y => m14_ns_1);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_0\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega16_2, B => CONFIG_rega9_0, C => 
        m18_0, D => un9_psel, Y => un271_psel);
    
    N_51_i : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PENABLE, B => 
        CoreAPB3_0_APBmslave0_PWRITE, C => \un30_psel\, D => 
        CoreAPB3_0_APBmslave7_PSELx, Y => N_51_i_0);
    
    \GEN_BITS.4.APB_32.un229_fixed_config\ : CFG2
      generic map(INIT => x"2")

      port map(A => \gpin2[4]_net_1\, B => \gpin3[4]_net_1\, Y
         => un229_fixed_config);
    
    g0_6_a3_0_4 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => g0_6_a3_0);
    
    \edge_both_RNO_0[10]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[10]_net_1\, B => N_65, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        \edge_both_RNO_0[10]_net_1\);
    
    \edge_both[0]\ : SLE
      port map(D => \edge_neg_7[0]\, CLK => FAB_CCC_GL0, EN => 
        edge_pos_2_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \edge_pos[0]\);
    
    \edge_pos_RNO[8]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[8]_net_1\, B => N_65, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        N_36_0);
    
    \GEN_BITS.27.APB_32.INTR_reg_277_ns_1[27]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_277_ns_1_1[27]\, B => 
        \CONFIG_reg_27[3]_net_1\, Y => \INTR_reg_277_ns_1[27]\);
    
    \CONFIG_reg_7[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un214_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_7[5]_net_1\);
    
    \CONFIG_reg_21[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un619_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_21[6]_net_1\);
    
    \gpin3[12]\ : SLE
      port map(D => \gpin2[12]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[12]_net_1\);
    
    \GEN_BITS.19.APB_32.edge_neg_197_iv_i_RNO[19]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[19]_net_1\, B => 
        \CONFIG_reg_19[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(19), Y => N_66_0);
    
    \GPOUT_reg_RNIMCCPA[5]\ : CFG4
      generic map(INIT => x"CC74")

      port map(A => m36_am_1, B => m36_ns_1_1, C => 
        \GPOUT_reg[5]_net_1\, D => m62_s_net_1, Y => m36_ns_1);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIQVH78\ : 
        CFG4
      generic map(INIT => x"2075")

      port map(A => m62_s_net_1, B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => \CONFIG_regrx[2]\, D
         => \GPOUT_reg_RNIQ6KF5[2]_net_1\, Y => m52_ns_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_12_RNI0M5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega20_2, B => CONFIG_rega12_1, C => 
        CONFIG_regro_12, D => CoreAPB3_0_APBmslave0_PADDR(6), Y
         => CONFIG_regria_12);
    
    \edge_both_RNO[20]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[20]\, B => \CONFIG_reg_20[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(20), Y => 
        \edge_neg_207[20]\);
    
    \INTR_reg[20]\ : SLE
      port map(D => \INTR_reg_207[20]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[20]_net_1\);
    
    \INTR_reg[13]\ : SLE
      port map(D => \INTR_reg_137[13]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[13]_net_1\);
    
    \edge_both_RNO_0[23]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_23[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_398_i_0);
    
    \INTR_reg_RNO_1[13]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_13[3]_net_1\, B => m161_ns_1, C
         => \edge_both[13]_net_1\, D => \CONFIG_reg_13[7]_net_1\, 
        Y => N_162_0);
    
    \INTR_reg_RNO_3[11]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_11[6]_net_1\, B => 
        \edge_pos[11]_net_1\, C => \gpin3[11]_net_1\, D => 
        \CONFIG_reg_11[7]_net_1\, Y => m146_ns_1);
    
    \GEN_BITS.29.APB_32.INTR_reg_297_ns_1[29]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_297_ns_1_1[29]\, B => 
        \CONFIG_reg_29[3]_net_1\, Y => \INTR_reg_297_ns_1[29]\);
    
    \edge_both[28]\ : SLE
      port map(D => \edge_neg_287[28]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_394_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[28]\);
    
    \GEN_BITS.17.APB_32.edge_both_177_iv_i[17]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[17]_net_1\, B => 
        \CONFIG_reg_17[3]_net_1\, C => un995_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(17), Y => 
        \edge_both_177_iv_i_0[17]\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_10\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \CONFIG_rega23_1\, B => CONFIG_rega3_0, C => 
        un9_psel, D => m18_0, Y => un98_psel);
    
    g0_2_0 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => g0_2_1_0);
    
    \GPOUT_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[7]_net_1\);
    
    \edge_both[29]\ : SLE
      port map(D => \edge_neg_297[29]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_396_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[29]\);
    
    \edge_both_RNO[21]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[21]\, B => \CONFIG_reg_21[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(21), Y => 
        \edge_neg_217[21]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_16\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un474_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_16);
    
    g0 : CFG4
      generic map(INIT => x"0020")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \g0_1\, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega1);
    
    \edge_neg[11]\ : SLE
      port map(D => \edge_neg_117_iv_i_0[11]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_436_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[11]_net_1\);
    
    \gpin1[10]\ : SLE
      port map(D => GPIO_IN_c(10), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[10]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0\ : 
        RAM64x18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => nc9, A_DOUT(7) => 
        \CONFIG_regrx[7]\, A_DOUT(6) => \CONFIG_regrx[6]\, 
        A_DOUT(5) => \CONFIG_regrx[5]\, A_DOUT(4) => 
        \CONFIG_regrx[4]\, A_DOUT(3) => \CONFIG_regrx[3]\, 
        A_DOUT(2) => \CONFIG_regrx[2]\, A_DOUT(1) => 
        \CONFIG_regrx[1]\, A_DOUT(0) => \CONFIG_regrx[0]\, 
        B_DOUT(17) => nc22, B_DOUT(16) => nc28, B_DOUT(15) => 
        nc14, B_DOUT(14) => nc5, B_DOUT(13) => nc21, B_DOUT(12)
         => nc15, B_DOUT(11) => nc3, B_DOUT(10) => nc10, 
        B_DOUT(9) => nc7, B_DOUT(8) => nc17, B_DOUT(7) => nc4, 
        B_DOUT(6) => nc12, B_DOUT(5) => nc2, B_DOUT(4) => nc23, 
        B_DOUT(3) => nc18, B_DOUT(2) => nc26, B_DOUT(1) => nc6, 
        B_DOUT(0) => nc11, BUSY => OPEN, A_ADDR_CLK => VCC_net_1, 
        A_DOUT_CLK => VCC_net_1, A_ADDR_SRST_N => VCC_net_1, 
        A_DOUT_SRST_N => VCC_net_1, A_ADDR_ARST_N => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_ADDR_EN => VCC_net_1, 
        A_DOUT_EN => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_ADDR(9) => GND_net_1, A_ADDR(8) => 
        GND_net_1, A_ADDR(7) => CoreAPB3_0_APBmslave0_PADDR(6), 
        A_ADDR(6) => CoreAPB3_0_APBmslave0_PADDR(5), A_ADDR(5)
         => CoreAPB3_0_APBmslave0_PADDR(4), A_ADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(3), A_ADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(2), A_ADDR(2) => GND_net_1, 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, 
        B_ADDR_CLK => VCC_net_1, B_DOUT_CLK => VCC_net_1, 
        B_ADDR_SRST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_ADDR_ARST_N => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, 
        B_ADDR_EN => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(1)
         => VCC_net_1, B_BLK(0) => VCC_net_1, B_ADDR(9) => 
        GND_net_1, B_ADDR(8) => GND_net_1, B_ADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(6), B_ADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(5), B_ADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(4), B_ADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(3), B_ADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(2), B_ADDR(2) => GND_net_1, 
        B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, C_CLK => 
        FAB_CCC_GL0, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => CoreAPB3_0_APBmslave0_PADDR(6), 
        C_ADDR(6) => CoreAPB3_0_APBmslave0_PADDR(5), C_ADDR(5)
         => CoreAPB3_0_APBmslave0_PADDR(4), C_ADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(3), C_ADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(2), C_ADDR(2) => GND_net_1, 
        C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, C_DIN(17)
         => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15) => 
        GND_net_1, C_DIN(14) => GND_net_1, C_DIN(13) => GND_net_1, 
        C_DIN(12) => GND_net_1, C_DIN(11) => GND_net_1, C_DIN(10)
         => GND_net_1, C_DIN(9) => GND_net_1, C_DIN(8) => 
        GND_net_1, C_DIN(7) => CoreAPB3_0_APBmslave0_PWDATA(7), 
        C_DIN(6) => CoreAPB3_0_APBmslave0_PWDATA(6), C_DIN(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), C_DIN(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), C_DIN(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), C_DIN(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), C_DIN(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), C_DIN(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), C_WEN => 
        CONFIG_reg_0_0_we, C_BLK(1) => VCC_net_1, C_BLK(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_ADDR_LAT => VCC_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => GND_net_1, 
        A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => VCC_net_1, B_EN
         => GND_net_1, B_ADDR_LAT => VCC_net_1, B_DOUT_LAT => 
        VCC_net_1, B_WIDTH(2) => GND_net_1, B_WIDTH(1) => 
        VCC_net_1, B_WIDTH(0) => VCC_net_1, C_EN => VCC_net_1, 
        C_WIDTH(2) => GND_net_1, C_WIDTH(1) => VCC_net_1, 
        C_WIDTH(0) => VCC_net_1, SII_LOCK => GND_net_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega6\ : CFG4
      generic map(INIT => x"0100")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => CONFIG_rega30_1, Y
         => CONFIG_rega6);
    
    \CONFIG_reg_30[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un880_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_30[6]_net_1\);
    
    \CONFIG_reg_28[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un822_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_28[7]_net_1\);
    
    \INTR_reg_RNO_1[16]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => \edge_pos[16]_net_1\, B => 
        \edge_neg[16]_net_1\, C => \CONFIG_reg_16[7]_net_1\, D
         => \CONFIG_reg_16[5]_net_1\, Y => 
        \INTR_reg_RNO_1[16]_net_1\);
    
    g0_10 : CFG4
      generic map(INIT => x"0020")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => g0_2_1_0, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega2);
    
    \GPOUT_reg[30]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(30), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_30);
    
    \INTR_reg[1]\ : SLE
      port map(D => N_6167_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[1]_net_1\);
    
    \edge_both[26]\ : SLE
      port map(D => \edge_neg_267[26]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_381_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[26]\);
    
    \INTR_reg_RNO_1[1]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_1[5]_net_1\, B => \edge_neg[1]\, 
        C => \CONFIG_reg_1[7]_net_1\, D => 
        \CONFIG_reg_1[6]_net_1\, Y => N_6177);
    
    \gpin2[14]\ : SLE
      port map(D => \gpin1[14]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[14]_net_1\);
    
    \edge_both_RNO_0[29]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_29[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_396_i_0);
    
    \CONFIG_reg_30[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un880_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_30[7]_net_1\);
    
    \INTR_reg[0]\ : SLE
      port map(D => N_6172_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[0]_net_1\);
    
    \edge_pos[15]\ : SLE
      port map(D => \edge_pos_157_iv_i_0[15]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_404_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[15]_net_1\);
    
    \GEN_BITS.15.APB_32.edge_pos_157_iv_i_RNO[15]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[15]_net_1\, B => 
        \CONFIG_reg_15[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(15), Y => N_198);
    
    \edge_pos_RNO_0[10]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[10]_net_1\, B => N_65, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        \edge_pos_RNO_0[10]_net_1\);
    
    \gpin1[18]\ : SLE
      port map(D => GPIO_IN_c(18), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[18]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_1\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un41_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_1);
    
    \CONFIG_reg_28[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un822_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_28[6]_net_1\);
    
    \CONFIG_reg_17[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un503_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_17[1]_net_1\);
    
    \edge_neg_RNO_0[10]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[10]_net_1\, B => N_65, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        \edge_neg_RNO_0[10]_net_1\);
    
    \CONFIG_reg_11_RNI84NL[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \gpin3[11]_net_1\, B => 
        \CONFIG_reg_11[1]_net_1\, Y => N_419_mux);
    
    m18 : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => m18_0, D => 
        CoreAPB3_0_APBmslave7_PSELx, Y => un11_psel_1_0);
    
    edge_neg_2_sqmuxa_428_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_14[3]_net_1\, D => un809_fixed_config, Y => 
        edge_neg_2_sqmuxa_428_i_0);
    
    \CONFIG_reg_11[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un329_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_11[1]_net_1\);
    
    \edge_both_RNO_0[26]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_26[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_381_i_0);
    
    \edge_both_RNO[12]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[12]_net_1\, B => N_296, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        i64_mux);
    
    \INTR_reg_RNING6H2[23]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[23]_net_1\, Y => INTR_reg_m_1);
    
    edge_pos_2_sqmuxa_387_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[7]_net_1\, B => N_65, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_387_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega18_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega18_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_25_RNI4N5U1\ : CFG3
      generic map(INIT => x"80")

      port map(A => CONFIG_rega25_2, B => CONFIG_regro_25, C => 
        CONFIG_rega25_0, Y => CONFIG_regria_25);
    
    edge_pos_2_sqmuxa_386_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_16[3]_net_1\, D => un901_fixed_config, Y => 
        edge_pos_2_sqmuxa_386_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_9_RNILMNR3\ : CFG4
      generic map(INIT => x"54FC")

      port map(A => g0_1_2, B => g0_i_a3_2_0, C => g0_i_a3_3_0, D
         => g0_i_0_1, Y => CONFIG_regror_23_1);
    
    \CONFIG_reg_1[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un41_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_1[3]_net_1\);
    
    \edge_both[13]\ : SLE
      port map(D => \edge_both_137_iv_i_0[13]\, CLK => 
        FAB_CCC_GL0, EN => N_211, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[13]_net_1\);
    
    \GEN_BITS.4.APB_32.un249_fixed_config\ : CFG2
      generic map(INIT => x"4")

      port map(A => \gpin2[4]_net_1\, B => \gpin3[4]_net_1\, Y
         => un249_fixed_config);
    
    \edge_pos_RNO_0[12]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[12]_net_1\, B => N_65, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        \edge_pos_RNO_0[12]_net_1\);
    
    \INTR_reg_RNO_3[15]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_15[6]_net_1\, B => 
        \edge_pos[15]_net_1\, C => \gpin3[15]_net_1\, D => 
        \CONFIG_reg_15[7]_net_1\, Y => m175_ns_1);
    
    \INTR_reg_RNO_2[8]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[8]_net_1\, B => 
        \CONFIG_reg_8[3]_net_1\, C => \edge_neg[8]_net_1\, D => 
        \CONFIG_reg_8[6]_net_1\, Y => N_6243);
    
    \GEN_BITS.22.APB_32.INTR_reg_227_ns_1_1[22]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_22[5]_net_1\, B => \edge_neg[22]\, 
        C => \CONFIG_reg_22[7]_net_1\, D => 
        \CONFIG_reg_22[6]_net_1\, Y => \INTR_reg_227_ns_1_1[22]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_31\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CONFIG_rega12_1, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un909_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_28\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un822_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_28);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_26_RNI5N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega26_1, B => CONFIG_rega26_2, C => 
        CONFIG_regro_26, D => CoreAPB3_0_APBmslave0_PADDR(4), Y
         => CONFIG_regria_26);
    
    edge_both_2_sqmuxa_452_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_11[3]_net_1\, D => un659_fixed_config, Y => 
        edge_both_2_sqmuxa_452_i_0);
    
    \INTR_reg_RNO_2[11]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[11]_net_1\, B => 
        \CONFIG_reg_11[3]_net_1\, C => \edge_neg[11]_net_1\, D
         => \CONFIG_reg_11[6]_net_1\, Y => N_150_0);
    
    \GPOUT_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[6]_net_1\);
    
    \CONFIG_reg_3[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un98_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_3[3]_net_1\);
    
    \GEN_BITS.13.APB_32.edge_neg_137_iv_i_RNO[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[13]_net_1\, B => 
        \CONFIG_reg_13[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(13), Y => N_186);
    
    \GEN_BITS.19.APB_32.un1107_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[19]_net_1\, B => \gpin3[19]_net_1\, Y
         => un1107_fixed_config);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_6\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega28_0, B => CONFIG_rega26_2, C => 
        m18_0, D => un9_psel, Y => un822_psel);
    
    \CONFIG_reg_2[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un69_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_2[6]_net_1\);
    
    \INTR_reg[31]\ : SLE
      port map(D => \INTR_reg_317[31]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[31]_net_1\);
    
    \GEN_BITS.18.APB_32.edge_neg_187_iv_i[18]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[18]_net_1\, B => N_101_0, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        \edge_neg_187_iv_i_0[18]\);
    
    \GEN_BITS.24.APB_32.INTR_reg_247_ns_1[24]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_247_ns_1_1[24]\, B => 
        \CONFIG_reg_24[3]_net_1\, Y => \INTR_reg_247_ns_1[24]\);
    
    \INTR_reg_RNO_0[10]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_10[7]_net_1\, B => 
        \CONFIG_reg_10[6]_net_1\, C => N_254, D => N_257, Y => 
        m259_ns_1);
    
    \gpin3[7]\ : SLE
      port map(D => \gpin2[7]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_20\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega2, Y
         => un69_psel);
    
    \GPOUT_reg_RNIQN3C5[11]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[11]_net_1\, B => 
        \INTR_reg[11]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => N_302);
    
    \GEN_BITS.22.APB_32.INTR_reg_227_ns_1[22]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_227_ns_1_1[22]\, B => 
        \CONFIG_reg_22[3]_net_1\, Y => \INTR_reg_227_ns_1[22]\);
    
    \edge_both_RNO[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[28]\, B => \CONFIG_reg_28[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(28), Y => 
        \edge_neg_287[28]\);
    
    edge_neg_2_sqmuxa_434_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_4[3]_net_1\, D => un249_fixed_config, Y => 
        edge_neg_2_sqmuxa_434_i_0);
    
    edge_both_2_sqmuxa_439_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_15[3]_net_1\, D => un883_fixed_config, Y => 
        edge_both_2_sqmuxa_439_i_0);
    
    edge_neg_2_sqmuxa_426_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_16[3]_net_1\, D => un921_fixed_config, Y => 
        edge_neg_2_sqmuxa_426_i_0);
    
    \GPOUT_reg[19]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(19), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[19]_net_1\);
    
    \GEN_BITS.26.APB_32.INTR_reg_267_ns_1_1[26]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_26[5]_net_1\, B => \edge_pos[26]\, 
        C => \CONFIG_reg_26[7]_net_1\, D => 
        \CONFIG_reg_26[6]_net_1\, Y => \INTR_reg_267_ns_1_1[26]\);
    
    \GEN_BITS.18.APB_32.edge_pos_187_iv_i_RNO[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[18]_net_1\, B => 
        \CONFIG_reg_18[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(18), Y => N_104_0);
    
    \GEN_BITS.13.APB_32.edge_both_137_iv_i_RNO[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[13]_net_1\, B => 
        \CONFIG_reg_13[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(13), Y => N_201);
    
    \gpin2[16]\ : SLE
      port map(D => \gpin1[16]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[16]_net_1\);
    
    \gpin2[9]\ : SLE
      port map(D => \gpin1[9]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[9]_net_1\);
    
    \edge_both_RNO_1[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[12]_net_1\, B => 
        \CONFIG_reg_12[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(12), Y => N_296);
    
    \edge_both[27]\ : SLE
      port map(D => \edge_neg_277[27]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_395_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[27]\);
    
    \CONFIG_reg_17_RNI2Q958[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_17[1]_net_1\, B => 
        \gpin3[17]_net_1\, C => \un3_prdata_o\, D => m332_ns_1, Y
         => N_333);
    
    \GEN_BITS.11.APB_32.edge_pos_117_iv_i[11]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[11]_net_1\, B => N_192, C => 
        \gpin3[11]_net_1\, D => \CONFIG_reg_11[3]_net_1\, Y => 
        \edge_pos_117_iv_i_0[11]\);
    
    \gpin3[11]\ : SLE
      port map(D => \gpin2[11]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[11]_net_1\);
    
    \INTR_reg_RNO[1]\ : CFG4
      generic map(INIT => x"DC10")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => N_65, C
         => \INTR_reg[1]_net_1\, D => \intr_3[1]\, Y => 
        N_6167_i_0);
    
    \CONFIG_reg_9[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un271_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_9[7]_net_1\);
    
    \GPOUT_reg[29]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(29), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_29);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_27\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un793_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_27);
    
    edge_pos_2_sqmuxa_404_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[15]_net_1\, B => N_65, C => 
        \gpin3[15]_net_1\, D => \CONFIG_reg_15[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_404_i_0);
    
    \GPOUT_reg_RNI66K552[5]\ : CFG4
      generic map(INIT => x"3373")

      port map(A => \CONFIG_regror_29\, B => m36_ns_1, C => 
        m62_s_net_1, D => \CONFIG_regror_28\, Y => N_37);
    
    m22_0_2 : CFG4
      generic map(INIT => x"0004")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \m22_0_2\);
    
    \INTR_reg_RNO_3[9]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => \edge_neg[9]_net_1\, B => \edge_pos[9]_net_1\, 
        C => \CONFIG_reg_9[6]_net_1\, D => 
        \CONFIG_reg_9[5]_net_1\, Y => m239_ns_1);
    
    \GEN_BITS.28.APB_32.INTR_reg_287_ns_1[28]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_287_ns_1_1[28]\, B => 
        \CONFIG_reg_28[3]_net_1\, Y => \INTR_reg_287_ns_1[28]\);
    
    \INTR_reg_RNO_1[0]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_0[5]_net_1\, B => \edge_pos[0]\, 
        C => \CONFIG_reg_0[7]_net_1\, D => 
        \CONFIG_reg_0[6]_net_1\, Y => m102_ns_1_0);
    
    \gpin2[6]\ : SLE
      port map(D => \gpin1[6]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[6]_net_1\);
    
    \gpin2[5]\ : SLE
      port map(D => \gpin1[5]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[5]_net_1\);
    
    \CONFIG_reg_9[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un271_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_9[1]_net_1\);
    
    g0_15 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega16_2);
    
    \GPOUT_reg_RNIUR3C5[13]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[13]_net_1\, B => 
        \INTR_reg[13]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => N_312);
    
    g0_0_1 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => \g0_0_1\);
    
    \edge_both[21]\ : SLE
      port map(D => \edge_neg_217[21]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_400_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[21]\);
    
    \INTR_reg_RNO_2[17]\ : CFG4
      generic map(INIT => x"5066")

      port map(A => \CONFIG_reg_17[5]_net_1\, B => 
        \gpin3[17]_net_1\, C => \edge_both[17]_net_1\, D => 
        \CONFIG_reg_17[7]_net_1\, Y => \INTR_reg_RNO_2[17]_net_1\);
    
    \INTR_reg[9]\ : SLE
      port map(D => \INTR_reg_97[9]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[9]_net_1\);
    
    \edge_neg_RNO_1[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[9]_net_1\, B => 
        \CONFIG_reg_9[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(9), Y => N_374);
    
    \CONFIG_reg_31[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un909_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_31[5]_net_1\);
    
    \gpin1[8]\ : SLE
      port map(D => GPIO_IN_c(8), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[8]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_24_RNIK9B11\ : CFG3
      generic map(INIT => x"80")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CONFIG_regro_24, C => CoreAPB3_0_APBmslave0_PADDR(5), Y
         => CONFIG_regria_24_0);
    
    \INTR_reg_RNO_2[15]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[15]_net_1\, B => 
        \CONFIG_reg_15[3]_net_1\, C => \edge_neg[15]_net_1\, D
         => \CONFIG_reg_15[6]_net_1\, Y => N_179);
    
    \edge_pos_RNO_1[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[9]_net_1\, B => 
        \CONFIG_reg_9[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(9), Y => N_377);
    
    \edge_both[22]\ : SLE
      port map(D => \edge_neg_227[22]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_392_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[22]\);
    
    \GPOUT_reg[31]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(31), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg_31\);
    
    \GEN_BITS.6.APB_32.edge_pos_67_iv_i_RNO[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[6]_net_1\, B => 
        \CONFIG_reg_6[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(6), Y => N_75_0);
    
    \CONFIG_reg_31[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un909_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_31[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_14\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega13, Y
         => un387_psel);
    
    \edge_pos_RNO[18]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[18]_net_1\, B => N_65, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        N_116_0);
    
    \CONFIG_reg_2[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un69_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_2[0]_net_1\);
    
    \INTR_reg[4]\ : SLE
      port map(D => \INTR_reg_47[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[4]_net_1\);
    
    \GPOUT_reg[8]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(8), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[8]_net_1\);
    
    \CONFIG_reg_5[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un156_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_5[5]_net_1\);
    
    \GEN_BITS.25.APB_32.INTR_reg_257_ns[25]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(25), B => N_65, 
        C => \INTR_reg[25]_net_1\, D => \INTR_reg_257_ns_1[25]\, 
        Y => \INTR_reg_257[25]\);
    
    \GPOUT_reg_RNIAKFJ5[4]\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \un30_psel\, B => m41_am_1, C => 
        \GPOUT_reg[4]_net_1\, Y => \GPOUT_reg_RNIAKFJ5[4]_net_1\);
    
    \INTR_reg_RNO_1[9]\ : CFG4
      generic map(INIT => x"D7DD")

      port map(A => \CONFIG_reg_9[3]_net_1\, B => m239_ns_1, C
         => \CONFIG_reg_9[6]_net_1\, D => \gpin3[9]_net_1\, Y => 
        N_240);
    
    \INTR_reg[19]\ : SLE
      port map(D => \INTR_reg_197[19]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[19]_net_1\);
    
    \GEN_BITS.18.APB_32.edge_both_187_iv_i[18]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[18]_net_1\, B => N_107_0, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        \edge_both_187_iv_i_0[18]\);
    
    \GEN_BITS.30.APB_32.INTR_reg_307_ns_1_1[30]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_30[5]_net_1\, B => \edge_neg[30]\, 
        C => \CONFIG_reg_30[7]_net_1\, D => 
        \CONFIG_reg_30[6]_net_1\, Y => \INTR_reg_307_ns_1_1[30]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega14_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega8_0);
    
    edge_both_2_sqmuxa_444_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_19[3]_net_1\, D => un1107_fixed_config, Y => 
        edge_both_2_sqmuxa_444_i_0);
    
    \GEN_BITS.19.APB_32.edge_pos_197_iv_i_RNO[19]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[19]_net_1\, B => 
        \CONFIG_reg_19[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(19), Y => N_72_0);
    
    \edge_neg[8]\ : SLE
      port map(D => \edge_neg_87_iv_i_0[8]\, CLK => FAB_CCC_GL0, 
        EN => N_37_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_neg[8]_net_1\);
    
    \edge_both[8]\ : SLE
      port map(D => \edge_both_87_iv_i_0[8]\, CLK => FAB_CCC_GL0, 
        EN => N_34_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_both[8]_net_1\);
    
    \INTR_reg_RNO_3[19]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_19[6]_net_1\, B => 
        \edge_pos[19]_net_1\, C => \gpin3[19]_net_1\, D => 
        \CONFIG_reg_19[7]_net_1\, Y => m58_1_ns_1);
    
    \CONFIG_reg_3[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un98_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_3[5]_net_1\);
    
    \edge_both[7]\ : SLE
      port map(D => \edge_both_77_iv_i_0[7]\, CLK => FAB_CCC_GL0, 
        EN => edge_both_2_sqmuxa_456_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[7]_net_1\);
    
    \CONFIG_reg_26[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un764_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_26[6]_net_1\);
    
    \GEN_BITS.14.APB_32.edge_neg_147_iv_i[14]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_neg[14]_net_1\, B => 
        \CONFIG_reg_14[3]_net_1\, C => un809_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(14), Y => 
        \edge_neg_147_iv_i_0[14]\);
    
    \CONFIG_reg_8[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un242_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_8[7]_net_1\);
    
    \CONFIG_reg_8[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un242_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_8[6]_net_1\);
    
    \CONFIG_reg_13_RNICCT7[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \gpin3[13]_net_1\, B => 
        \CONFIG_reg_13[1]_net_1\, Y => N_421_mux);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega30_1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega30_1);
    
    \CONFIG_reg_14[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un416_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_14[7]_net_1\);
    
    \gpin3[13]\ : SLE
      port map(D => \gpin2[13]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[13]_net_1\);
    
    \CONFIG_reg_6[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un185_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_6[3]_net_1\);
    
    m24 : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \m22_0_2\, D => 
        un1_psel_280_2, Y => \un3_prdata_o\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega5_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega5_0);
    
    \edge_neg[10]\ : SLE
      port map(D => N_48, CLK => FAB_CCC_GL0, EN => 
        \edge_neg_RNO_0[10]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[10]_net_1\);
    
    \GEN_BITS.14.APB_32.un809_fixed_config\ : CFG2
      generic map(INIT => x"4")

      port map(A => \gpin2[14]_net_1\, B => \gpin3[14]_net_1\, Y
         => un809_fixed_config);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_12\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un358_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_12);
    
    \CONFIG_reg_24[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un706_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_24[3]_net_1\);
    
    \INTR_reg_RNO_3[7]\ : CFG3
      generic map(INIT => x"35")

      port map(A => \edge_pos[7]_net_1\, B => \edge_neg[7]_net_1\, 
        C => \CONFIG_reg_7[5]_net_1\, Y => N_6193);
    
    \INTR_reg[3]\ : SLE
      port map(D => N_6165_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[3]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_26\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un764_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_26);
    
    \INTR_reg_RNO_0[11]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_11[7]_net_1\, B => 
        \CONFIG_reg_11[5]_net_1\, C => N_147_0, D => N_150_0, Y
         => m152_ns_1);
    
    \GEN_BITS.14.APB_32.un789_fixed_config\ : CFG2
      generic map(INIT => x"2")

      port map(A => \gpin2[14]_net_1\, B => \gpin3[14]_net_1\, Y
         => un789_fixed_config);
    
    \INTR_reg_RNO_1[10]\ : CFG4
      generic map(INIT => x"8882")

      port map(A => \CONFIG_reg_10[3]_net_1\, B => m253_ns_1_0, C
         => \CONFIG_reg_10[7]_net_1\, D => \gpin3[10]_net_1\, Y
         => N_254);
    
    \edge_both[25]\ : SLE
      port map(D => \edge_neg_257[25]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_382_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[25]\);
    
    \CONFIG_reg_1[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un41_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_1[6]_net_1\);
    
    edge_both_2_sqmuxa_458_i : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[5]_net_1\, B => N_65, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        edge_both_2_sqmuxa_458_i_0);
    
    \CONFIG_reg_23[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un677_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_23[3]_net_1\);
    
    m23_0 : CFG3
      generic map(INIT => x"20")

      port map(A => \m22_0_2\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => un1_psel_280_2, Y
         => \N_6186\);
    
    \INTR_reg_RNO[2]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[2]_net_1\, B => N_6195, C => 
        CoreAPB3_0_APBmslave0_PWDATA(2), D => N_65, Y => 
        N_6196_i_0);
    
    \INTR_reg_RNO_1[8]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_8[3]_net_1\, B => m14_ns_1, C => 
        \edge_both[8]_net_1\, D => \CONFIG_reg_8[7]_net_1\, Y => 
        N_15_0);
    
    \CONFIG_reg_7[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un214_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_7[1]_net_1\);
    
    \INTR_reg_RNIPI6H2[25]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[25]_net_1\, Y => N_435);
    
    \GPOUT_reg[9]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(9), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[9]_net_1\);
    
    g0_3 : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega21_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_2\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un69_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_2);
    
    \CONFIG_reg_9_RNI1T7S7[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_9[1]_net_1\, B => 
        \gpin3[9]_net_1\, C => \un3_prdata_o\, D => m352_ns_1, Y
         => N_353);
    
    \GEN_BITS.29.APB_32.INTR_reg_297_ns_1_1[29]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_29[5]_net_1\, B => \edge_neg[29]\, 
        C => \CONFIG_reg_29[7]_net_1\, D => 
        \CONFIG_reg_29[6]_net_1\, Y => \INTR_reg_297_ns_1_1[29]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_3_RNIGVHT1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega0_2, B => \CONFIG_rega23_1\, C => 
        CONFIG_regro_3, D => CoreAPB3_0_APBmslave0_PADDR(6), Y
         => CONFIG_regria_3);
    
    g0_i_a3_0 : CFG2
      generic map(INIT => x"7")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => g0_i_a3_2_0);
    
    \GEN_BITS.29.APB_32.INTR_reg_297_ns[29]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(29), B => N_65, 
        C => \INTR_reg[29]_net_1\, D => \INTR_reg_297_ns_1[29]\, 
        Y => \INTR_reg_297[29]\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_24\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega20, Y
         => un590_psel);
    
    \INTR_reg_RNO_1[3]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_3[5]_net_1\, B => \edge_neg[3]\, 
        C => \CONFIG_reg_3[7]_net_1\, D => 
        \CONFIG_reg_3[6]_net_1\, Y => N_6174);
    
    \INTR_reg_RNO[7]\ : CFG4
      generic map(INIT => x"330A")

      port map(A => \INTR_reg[7]_net_1\, B => N_6158, C => 
        CoreAPB3_0_APBmslave0_PWDATA(7), D => N_65, Y => 
        N_6160_i_0);
    
    \CONFIG_reg_31[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un909_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_31[6]_net_1\);
    
    \gpin1[12]\ : SLE
      port map(D => GPIO_IN_c(12), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[12]_net_1\);
    
    \GEN_BITS.26.APB_32.INTR_reg_267_ns[26]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(26), B => N_65, 
        C => \INTR_reg[26]_net_1\, D => \INTR_reg_267_ns_1[26]\, 
        Y => \INTR_reg_267[26]\);
    
    \edge_both[18]\ : SLE
      port map(D => \edge_both_187_iv_i_0[18]\, CLK => 
        FAB_CCC_GL0, EN => N_115_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[18]_net_1\);
    
    \GEN_BITS.28.APB_32.INTR_reg_287_ns_1_1[28]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_28[5]_net_1\, B => \edge_neg[28]\, 
        C => \CONFIG_reg_28[7]_net_1\, D => 
        \CONFIG_reg_28[6]_net_1\, Y => \INTR_reg_287_ns_1_1[28]\);
    
    edge_neg_2_sqmuxa_423_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[19]_net_1\, B => N_65, C => 
        \gpin3[19]_net_1\, D => \CONFIG_reg_19[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_423_i_0);
    
    \CONFIG_reg_13[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un387_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_13[1]_net_1\);
    
    \INTR_reg[12]\ : SLE
      port map(D => \INTR_reg_127[12]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[12]_net_1\);
    
    \edge_both[19]\ : SLE
      port map(D => \edge_both_197_iv_i_0[19]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_444_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[19]_net_1\);
    
    edge_both_2_sqmuxa_456_i : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[7]_net_1\, B => N_65, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        edge_both_2_sqmuxa_456_i_0);
    
    m26 : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => \m22_0_2\, D => 
        CONFIG_rega11_2, Y => \un30_psel\);
    
    \GEN_BITS.7.APB_32.edge_both_77_iv_i_RNO[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[7]_net_1\, B => 
        \CONFIG_reg_7[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(7), Y => N_6190);
    
    \edge_both[4]\ : SLE
      port map(D => \edge_both_47_iv_i_0[4]\, CLK => FAB_CCC_GL0, 
        EN => edge_both_2_sqmuxa_446_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[4]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIADDB8\ : 
        CFG4
      generic map(INIT => x"4073")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        m62_s_net_1, C => \CONFIG_regrx[4]\, D => 
        \GPOUT_reg_RNIAKFJ5[4]_net_1\, Y => N_92_i_1_1);
    
    g0_5_0_a3 : CFG4
      generic map(INIT => x"0040")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \g0_5_0_a3_1\, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega4);
    
    \GEN_BITS.5.APB_32.edge_both_57_iv_i_RNO[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[5]_net_1\, B => 
        \CONFIG_reg_5[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(5), Y => N_6152);
    
    \GEN_BITS.19.APB_32.edge_both_197_iv_i[19]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[19]_net_1\, B => 
        \CONFIG_reg_19[3]_net_1\, C => un1107_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(19), Y => 
        \edge_both_197_iv_i_0[19]\);
    
    \edge_neg_RNO_0[12]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[12]_net_1\, B => N_65, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        \edge_neg_RNO_0[12]_net_1\);
    
    \edge_neg_RNO[9]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[9]_net_1\, B => N_374, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        N_460_mux);
    
    \INTR_reg_RNO_2[19]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[19]_net_1\, B => 
        \CONFIG_reg_19[3]_net_1\, C => \edge_neg[19]_net_1\, D
         => \CONFIG_reg_19[6]_net_1\, Y => N_62_0);
    
    \GEN_BITS.21.APB_32.INTR_reg_217_ns[21]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(21), B => N_65, 
        C => \INTR_reg[21]_net_1\, D => \INTR_reg_217_ns_1[21]\, 
        Y => \INTR_reg_217[21]\);
    
    \CONFIG_reg_15[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un445_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_15[3]_net_1\);
    
    \GEN_BITS.31.APB_32.INTR_reg_317_ns_1[31]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_317_ns_1_1[31]\, B => 
        \CONFIG_reg_31[3]_net_1\, Y => \INTR_reg_317_ns_1[31]\);
    
    \CONFIG_reg_5[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un156_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_5[1]_net_1\);
    
    \edge_neg[13]\ : SLE
      port map(D => \edge_neg_137_iv_i_0[13]\, CLK => FAB_CCC_GL0, 
        EN => N_215, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_neg[13]_net_1\);
    
    \INTR_reg_RNO_0[17]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \CONFIG_reg_17[6]_net_1\, B => 
        \CONFIG_reg_17[3]_net_1\, C => \INTR_reg_RNO_1[17]_net_1\, 
        D => \INTR_reg_RNO_2[17]_net_1\, Y => N_126_0);
    
    \edge_both[16]\ : SLE
      port map(D => \edge_both_167_iv_i_0[16]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_462_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[16]_net_1\);
    
    \GEN_BITS.4.REG_INT.intr_9_u_ns_1[4]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \edge_both[4]_net_1\, B => 
        \CONFIG_reg_4[6]_net_1\, C => \CONFIG_reg_4[5]_net_1\, Y
         => \intr_9_u_ns_1[4]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_4\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un127_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_4);
    
    \GEN_BITS.4.APB_32.un267_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[4]_net_1\, B => \gpin3[4]_net_1\, Y
         => un267_fixed_config);
    
    \CONFIG_reg_12[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un358_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_12[6]_net_1\);
    
    \m62_s\ : CFG4
      generic map(INIT => x"8FFF")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \m22_0_2\, D => 
        un1_psel_280_2, Y => m62_s_net_1);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_27_RNI6N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega30_2, B => \CONFIG_rega23_1\, C
         => CONFIG_regro_27, D => CoreAPB3_0_APBmslave0_PADDR(4), 
        Y => CONFIG_regria_27);
    
    \CONFIG_reg_14[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un416_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_14[6]_net_1\);
    
    \gpin2[17]\ : SLE
      port map(D => \gpin1[17]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[17]_net_1\);
    
    \edge_pos[19]\ : SLE
      port map(D => \edge_pos_197_iv_i_0[19]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_402_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[19]_net_1\);
    
    \GPOUT_reg_RNISP3C5[12]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[12]_net_1\, B => 
        \INTR_reg[12]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => m309_ns_1);
    
    \CONFIG_reg_10[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un300_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_10[3]_net_1\);
    
    \INTR_reg_RNO_0[15]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_15[7]_net_1\, B => 
        \CONFIG_reg_15[5]_net_1\, C => N_176, D => N_179, Y => 
        m181_ns_1);
    
    \INTR_reg[16]\ : SLE
      port map(D => \INTR_reg_167[16]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[16]_net_1\);
    
    \GPOUT_reg_RNI6JKF5[8]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[8]_net_1\, B => 
        \INTR_reg[8]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => N_345);
    
    \gpin1[9]\ : SLE
      port map(D => GPIO_IN_c(9), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[9]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_15\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un445_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_15);
    
    \GEN_BITS.28.APB_32.INTR_reg_287_ns[28]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(28), B => N_65, 
        C => \INTR_reg[28]_net_1\, D => \INTR_reg_287_ns_1[28]\, 
        Y => \INTR_reg_287[28]\);
    
    \CONFIG_reg_19[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un561_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_19[5]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_9_RNIC1BA1\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CONFIG_regro_9, C => CoreAPB3_0_APBmslave0_PADDR(6), D
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => g0_i_a3_3_0);
    
    \edge_both_RNO_0[3]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_3[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_377_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_11\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un329_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_11);
    
    \CONFIG_reg_13[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un387_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_13[7]_net_1\);
    
    \GPOUT_reg_RNIA84C5[19]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[19]_net_1\, B => 
        \INTR_reg[19]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => m342_ns_1);
    
    \GEN_BITS.5.APB_32.edge_pos_57_iv_i[5]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[5]_net_1\, B => N_70, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        \edge_pos_57_iv_i_0[5]\);
    
    \gpin2[7]\ : SLE
      port map(D => \gpin1[7]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_19\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega17, Y
         => un503_psel);
    
    \GPOUT_reg_RNITGG25[15]\ : CFG4
      generic map(INIT => x"15BF")

      port map(A => \N_6186\, B => \un30_psel\, C => 
        \GPOUT_reg[15]_net_1\, D => \INTR_reg[15]_net_1\, Y => 
        m323_ns_1);
    
    \INTR_reg_RNO[8]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[8]_net_1\, B => m20_0_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(8), D => N_65, Y => 
        \INTR_reg_87[8]\);
    
    \GPOUT_reg[10]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(10), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[10]_net_1\);
    
    \GPOUT_reg_RNI644C5[17]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[17]_net_1\, B => 
        \INTR_reg[17]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => m332_ns_1);
    
    \CONFIG_reg_26[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un764_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_26[3]_net_1\);
    
    \edge_neg[9]\ : SLE
      port map(D => N_460_mux, CLK => FAB_CCC_GL0, EN => N_381, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \edge_neg[9]_net_1\);
    
    \gpin3[5]\ : SLE
      port map(D => \gpin2[5]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[5]_net_1\);
    
    \GEN_BITS.18.APB_32.edge_both_187_iv_i_RNO[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[18]_net_1\, B => 
        \CONFIG_reg_18[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(18), Y => N_107_0);
    
    \GEN_BITS.7.APB_32.edge_neg_77_iv_i[7]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[7]_net_1\, B => N_6192, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        \edge_neg_77_iv_i_0[7]\);
    
    \CONFIG_reg_29[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un851_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_29[3]_net_1\);
    
    \GPOUT_reg[13]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(13), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[13]_net_1\);
    
    \gpin3[6]\ : SLE
      port map(D => \gpin2[6]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[6]_net_1\);
    
    \edge_neg[5]\ : SLE
      port map(D => \edge_neg_57_iv_i_0[5]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_410_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[5]_net_1\);
    
    \CONFIG_reg_15[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un445_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_15[1]_net_1\);
    
    \CONFIG_reg_3[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un98_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_3[6]_net_1\);
    
    \CONFIG_reg_23[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un677_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_23[5]_net_1\);
    
    \CONFIG_reg_18[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un532_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_18[3]_net_1\);
    
    g0_12 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega0_2);
    
    \GPOUT_reg[20]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(20), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_20);
    
    m18_0_0 : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => m18_0);
    
    \edge_both[3]\ : SLE
      port map(D => \edge_neg_37[3]\, CLK => FAB_CCC_GL0, EN => 
        edge_pos_2_sqmuxa_377_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[3]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_7\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un214_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_7);
    
    \INTR_reg[7]\ : SLE
      port map(D => N_6160_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[7]_net_1\);
    
    m7_0 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), Y => un1_psel_280_2);
    
    \gpin2[15]\ : SLE
      port map(D => \gpin1[15]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[15]_net_1\);
    
    \GPOUT_reg[23]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(23), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_23);
    
    \INTR_reg_RNO_0[9]\ : CFG3
      generic map(INIT => x"2E")

      port map(A => N_240, B => \CONFIG_reg_9[7]_net_1\, C => 
        N_433_mux, Y => m244_ns_1);
    
    \GPOUT_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[1]_net_1\);
    
    \GEN_BITS.8.APB_32.edge_neg_87_iv_i_RNO[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[8]_net_1\, B => 
        \CONFIG_reg_8[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(8), Y => N_22_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_0\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un11_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_9\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un271_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_9);
    
    \CONFIG_reg_19[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un561_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_19[6]_net_1\);
    
    \GEN_BITS.4.REG_INT.intr_9_u_bm[4]\ : CFG4
      generic map(INIT => x"BE14")

      port map(A => \CONFIG_reg_4[6]_net_1\, B => 
        \CONFIG_reg_4[5]_net_1\, C => \gpin3[4]_net_1\, D => 
        N_5144, Y => \intr_9_u_bm[4]\);
    
    \gpin3[14]\ : SLE
      port map(D => \gpin2[14]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[14]_net_1\);
    
    \INTR_reg_RNO_1[11]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_11[3]_net_1\, B => m146_ns_1, C
         => \edge_both[11]_net_1\, D => \CONFIG_reg_11[7]_net_1\, 
        Y => N_147_0);
    
    \CONFIG_reg_20[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un590_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_20[5]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_11\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega25_2, B => CONFIG_rega25_0, C => 
        un9_psel, D => m18_0, Y => un735_psel);
    
    \GEN_BITS.27.APB_32.INTR_reg_277_ns_1_1[27]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_27[5]_net_1\, B => \edge_neg[27]\, 
        C => \CONFIG_reg_27[7]_net_1\, D => 
        \CONFIG_reg_27[6]_net_1\, Y => \INTR_reg_277_ns_1_1[27]\);
    
    \GEN_BITS.25.APB_32.INTR_reg_257_ns_1_1[25]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_25[5]_net_1\, B => \edge_neg[25]\, 
        C => \CONFIG_reg_25[7]_net_1\, D => 
        \CONFIG_reg_25[6]_net_1\, Y => \INTR_reg_257_ns_1_1[25]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_27\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CONFIG_rega30_2, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un793_psel);
    
    \edge_both_RNO_0[0]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_0[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_i_0);
    
    \GEN_BITS.6.APB_32.edge_both_67_iv_i[6]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[6]_net_1\, B => 
        \CONFIG_reg_6[3]_net_1\, C => un379_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(6), Y => 
        \edge_both_67_iv_i_0[6]\);
    
    \CONFIG_reg_7[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un214_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_7[6]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_13\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega18, Y
         => un532_psel);
    
    \edge_both[1]\ : SLE
      port map(D => \edge_neg_17[1]\, CLK => FAB_CCC_GL0, EN => 
        edge_pos_2_sqmuxa_399_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[1]\);
    
    \edge_pos[14]\ : SLE
      port map(D => \edge_pos_147_iv_i_0[14]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_379_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[14]_net_1\);
    
    \GEN_BITS.2.REG_GPOUT.GPIO_OUT_i_5[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG_reg_2[0]_net_1\, B => 
        \GPOUT_reg[2]_net_1\, Y => GPIO_OUT_c(2));
    
    \edge_both[17]\ : SLE
      port map(D => \edge_both_177_iv_i_0[17]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_437_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[17]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_29_RNI8N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega21_1, B => CONFIG_rega30_2, C => 
        CONFIG_regro_29, D => CoreAPB3_0_APBmslave0_PADDR(3), Y
         => CONFIG_regria_29);
    
    \INTR_reg_RNO_0[8]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_8[7]_net_1\, B => 
        \CONFIG_reg_8[5]_net_1\, C => N_15_0, D => N_6243, Y => 
        m20_0_ns_1);
    
    edge_neg_2_sqmuxa_427_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[15]_net_1\, B => N_65, C => 
        \gpin3[15]_net_1\, D => \CONFIG_reg_15[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_427_i_0);
    
    \edge_both_RNO[27]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[27]\, B => \CONFIG_reg_27[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(27), Y => 
        \edge_neg_277[27]\);
    
    \INTR_reg[21]\ : SLE
      port map(D => \INTR_reg_217[21]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[21]_net_1\);
    
    \GEN_BITS.20.APB_32.INTR_reg_207_ns_1_1[20]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_20[5]_net_1\, B => \edge_neg[20]\, 
        C => \CONFIG_reg_20[7]_net_1\, D => 
        \CONFIG_reg_20[6]_net_1\, Y => \INTR_reg_207_ns_1_1[20]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega25_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega25_2);
    
    \GEN_BITS.7.APB_32.edge_both_77_iv_i[7]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[7]_net_1\, B => N_6190, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        \edge_both_77_iv_i_0[7]\);
    
    \edge_both_RNO_0[24]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_24[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_397_i_0);
    
    \GEN_BITS.0.REG_GEN.un9_psel\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_48_1, B => m46_1_0, C => 
        CoreAPB3_0_APBmslave0_PWRITE, D => 
        CoreAPB3_0_APBmslave0_PENABLE, Y => un9_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_5_RNILMNR3\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => CONFIG_regria_24_0, B => CONFIG_regria_5_0, C
         => CONFIG_rega5_0, D => CONFIG_rega24_0, Y => 
        CONFIG_regror_2);
    
    \gpin1[11]\ : SLE
      port map(D => GPIO_IN_c(11), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[11]_net_1\);
    
    \edge_both_RNO_1[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[9]_net_1\, B => 
        \CONFIG_reg_9[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(9), Y => N_288);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_30_RNI0O5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega30_1, B => CONFIG_rega30_2, C => 
        CONFIG_regro_30, D => CoreAPB3_0_APBmslave0_PADDR(2), Y
         => CONFIG_regria_30);
    
    \edge_neg[7]\ : SLE
      port map(D => \edge_neg_77_iv_i_0[7]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_408_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[7]_net_1\);
    
    \INTR_reg_RNILF7H2[30]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[30]_net_1\, Y => N_439);
    
    \edge_both[11]\ : SLE
      port map(D => \edge_both_117_iv_i_0[11]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_452_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[11]_net_1\);
    
    \GEN_BITS.31.REG_GPOUT.GPIO_OUT_i_63[31]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG_reg_31[0]_net_1\, B => \GPOUT_reg_31\, 
        Y => USB_RST_c);
    
    \GEN_BITS.15.APB_32.edge_pos_157_iv_i[15]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[15]_net_1\, B => N_198, C => 
        \gpin3[15]_net_1\, D => \CONFIG_reg_15[3]_net_1\, Y => 
        \edge_pos_157_iv_i_0[15]\);
    
    \CONFIG_reg_15_RNILUFP7[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_15[1]_net_1\, B => 
        \gpin3[15]_net_1\, C => \un3_prdata_o\, D => m323_ns_1, Y
         => N_324);
    
    \INTR_reg_RNO_0[19]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \CONFIG_reg_19[7]_net_1\, B => 
        \CONFIG_reg_19[5]_net_1\, C => N_59_0, D => N_62_0, Y => 
        m64_1_ns_1);
    
    \GEN_BITS.24.APB_32.INTR_reg_247_ns_1_1[24]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_24[5]_net_1\, B => \edge_neg[24]\, 
        C => \CONFIG_reg_24[7]_net_1\, D => 
        \CONFIG_reg_24[6]_net_1\, Y => \INTR_reg_247_ns_1_1[24]\);
    
    \INTR_reg[2]\ : SLE
      port map(D => N_6196_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[2]_net_1\);
    
    \INTR_reg_RNO_1[17]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => \edge_pos[17]_net_1\, B => 
        \edge_neg[17]_net_1\, C => \CONFIG_reg_17[7]_net_1\, D
         => \CONFIG_reg_17[5]_net_1\, Y => 
        \INTR_reg_RNO_1[17]_net_1\);
    
    \edge_both[12]\ : SLE
      port map(D => i64_mux, CLK => FAB_CCC_GL0, EN => 
        \edge_both_RNO_0[12]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[12]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_19\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un561_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_19);
    
    \GEN_BITS.19.APB_32.edge_pos_197_iv_i[19]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[19]_net_1\, B => N_72_0, C => 
        \gpin3[19]_net_1\, D => \CONFIG_reg_19[3]_net_1\, Y => 
        \edge_pos_197_iv_i_0[19]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_19\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CONFIG_rega0_2, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un561_psel);
    
    \GEN_BITS.11.APB_32.edge_pos_117_iv_i_RNO[11]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[11]_net_1\, B => 
        \CONFIG_reg_11[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(11), Y => N_192);
    
    \CONFIG_reg_9[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un271_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_9[5]_net_1\);
    
    \edge_neg[14]\ : SLE
      port map(D => \edge_neg_147_iv_i_0[14]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_428_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[14]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_0_RNIUNO0P\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => CONFIG_regror_17, B => CONFIG_regror_19, C
         => CONFIG_regror_18, D => CONFIG_regror_16, Y => 
        \CONFIG_regror_28\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega26_2, B => CONFIG_rega16_0, C => 
        un9_psel, D => m18_0, Y => un474_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_22\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un648_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_22);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_6_RNI7V3R3\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => CONFIG_regro_6, B => CONFIG_regro_7, C => 
        CONFIG_rega7, D => CONFIG_rega6, Y => CONFIG_regror_11);
    
    \edge_pos[18]\ : SLE
      port map(D => \edge_pos_187_iv_i_0[18]\, CLK => FAB_CCC_GL0, 
        EN => N_116_0, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_pos[18]_net_1\);
    
    \edge_pos_RNO_0[9]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[9]_net_1\, B => N_65, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        N_382);
    
    \INTR_reg_RNO_1[15]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_15[3]_net_1\, B => m175_ns_1, C
         => \edge_both[15]_net_1\, D => \CONFIG_reg_15[7]_net_1\, 
        Y => N_176);
    
    \INTR_reg_RNIKD6H2[20]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[20]_net_1\, Y => N_438);
    
    \edge_both[6]\ : SLE
      port map(D => \edge_both_67_iv_i_0[6]\, CLK => FAB_CCC_GL0, 
        EN => edge_both_2_sqmuxa_457_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[6]_net_1\);
    
    \GEN_BITS.8.APB_32.edge_neg_87_iv_i[8]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[8]_net_1\, B => N_22_0, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        \edge_neg_87_iv_i_0[8]\);
    
    \edge_both[20]\ : SLE
      port map(D => \edge_neg_207[20]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_401_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[20]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_23_RNIGRQJB\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => CONFIG_regror_23_1, B => CONFIG_regria_25, C
         => CONFIG_regria_23, D => CONFIG_regror_2, Y => 
        CONFIG_regror_23);
    
    \INTR_reg[10]\ : SLE
      port map(D => \INTR_reg_107[10]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[10]_net_1\);
    
    \GEN_BITS.7.APB_32.edge_pos_77_iv_i_RNO[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[7]_net_1\, B => 
        \CONFIG_reg_7[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(7), Y => N_6191);
    
    \CONFIG_reg_18[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un532_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_18[1]_net_1\);
    
    \GPOUT_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[5]_net_1\);
    
    \gpin3[16]\ : SLE
      port map(D => \gpin2[16]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[16]_net_1\);
    
    \INTR_reg_RNO_0[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => m67_0_ns_1_0, B => \CONFIG_reg_2[3]_net_1\, Y
         => N_6195);
    
    \GEN_BITS.17.APB_32.edge_pos_177_iv_i[17]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_pos[17]_net_1\, B => 
        \CONFIG_reg_17[3]_net_1\, C => un957_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(17), Y => 
        \edge_pos_177_iv_i_0[17]\);
    
    \edge_both_RNO[13]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[13]_net_1\, B => N_65, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        N_211);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_21\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega1, Y
         => un41_psel);
    
    \CONFIG_reg_4[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un127_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_4[6]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_11\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CONFIG_rega11_2, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un329_psel);
    
    \INTR_reg_RNO_0[5]\ : CFG4
      generic map(INIT => x"5702")

      port map(A => \CONFIG_reg_5[6]_net_1\, B => 
        \CONFIG_reg_5[7]_net_1\, C => N_88, D => N_6163, Y => 
        N_90);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_16_RNI4M5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega16_2, B => CONFIG_rega26_2, C => 
        CONFIG_regro_16, D => CoreAPB3_0_APBmslave0_PADDR(5), Y
         => CONFIG_regria_16);
    
    \GPOUT_reg[11]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(11), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[11]_net_1\);
    
    \edge_neg_RNO[13]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[13]_net_1\, B => N_65, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        N_215);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega26_2, B => CONFIG_rega22_0, C => 
        un9_psel, D => m18_0, Y => un648_psel);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_23\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega26, Y
         => un764_psel);
    
    \edge_both_RNO_0[20]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_20[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_401_i_0);
    
    \GEN_BITS.19.APB_32.edge_neg_197_iv_i[19]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[19]_net_1\, B => N_66_0, C => 
        \gpin3[19]_net_1\, D => \CONFIG_reg_19[3]_net_1\, Y => 
        \edge_neg_197_iv_i_0[19]\);
    
    \edge_pos[10]\ : SLE
      port map(D => N_44, CLK => FAB_CCC_GL0, EN => 
        \edge_pos_RNO_0[10]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[10]_net_1\);
    
    \gpin2[19]\ : SLE
      port map(D => \gpin1[19]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[19]_net_1\);
    
    \edge_neg_RNO_0[9]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[9]_net_1\, B => N_65, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        N_381);
    
    \INTR_reg[6]\ : SLE
      port map(D => \INTR_reg_67[6]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[6]_net_1\);
    
    edge_pos_2_sqmuxa_383_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[11]_net_1\, B => N_65, C => 
        \gpin3[11]_net_1\, D => \CONFIG_reg_11[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_383_i_0);
    
    \GPOUT_reg[17]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(17), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[17]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_6\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un185_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_6);
    
    \edge_both_RNO[22]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[22]\, B => \CONFIG_reg_22[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(22), Y => 
        \edge_neg_227[22]\);
    
    \INTR_reg_RNIOH6H2[24]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[24]_net_1\, Y => N_436);
    
    \CONFIG_reg_7_RNIRN803[1]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => \INTR_reg[7]_net_1\, B => 
        \CONFIG_reg_7[1]_net_1\, C => \un3_prdata_o\, D => 
        \gpin3[7]_net_1\, Y => m23_am_1);
    
    \GPOUT_reg[21]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(21), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_21);
    
    \INTR_reg_RNO_2[14]\ : CFG4
      generic map(INIT => x"5066")

      port map(A => \CONFIG_reg_14[5]_net_1\, B => 
        \gpin3[14]_net_1\, C => \edge_both[14]_net_1\, D => 
        \CONFIG_reg_14[7]_net_1\, Y => \INTR_reg_RNO_2[14]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_15\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega10, Y
         => un300_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_17_RNII0AC2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => 
        CONFIG_regrff_17_RNI3JFF1, Y => CONFIG_regror_10);
    
    \GPOUT_reg[27]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(27), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_27);
    
    g0_1 : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => g0_1_2, Y => 
        CONFIG_rega20);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_21_RNI0N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega21_1, B => CONFIG_rega25_2, C => 
        CONFIG_regro_21, D => CoreAPB3_0_APBmslave0_PADDR(5), Y
         => CONFIG_regria_21);
    
    \gpin1[13]\ : SLE
      port map(D => GPIO_IN_c(13), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[13]_net_1\);
    
    \GEN_BITS.5.APB_32.edge_neg_57_iv_i[5]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[5]_net_1\, B => N_6155, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        \edge_neg_57_iv_i_0[5]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega29_0\ : CFG3
      generic map(INIT => x"20")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => CONFIG_rega29_0);
    
    \edge_neg[16]\ : SLE
      port map(D => \edge_neg_167_iv_i_0[16]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_426_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[16]_net_1\);
    
    \CONFIG_reg_4[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un127_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_4[3]_net_1\);
    
    edge_both_2_sqmuxa_457_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_6[3]_net_1\, D => un379_fixed_config, Y => 
        edge_both_2_sqmuxa_457_i_0);
    
    \edge_both[15]\ : SLE
      port map(D => \edge_both_157_iv_i_0[15]\, CLK => 
        FAB_CCC_GL0, EN => edge_both_2_sqmuxa_439_i_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \edge_both[15]_net_1\);
    
    edge_pos_2_sqmuxa_390_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_17[3]_net_1\, D => un957_fixed_config, Y => 
        edge_pos_2_sqmuxa_390_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_3\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un98_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_3);
    
    \GEN_BITS.15.APB_32.edge_neg_157_iv_i[15]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[15]_net_1\, B => N_189, C => 
        \gpin3[15]_net_1\, D => \CONFIG_reg_15[3]_net_1\, Y => 
        \edge_neg_157_iv_i_0[15]\);
    
    \GEN_BITS.14.APB_32.edge_pos_147_iv_i[14]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_pos[14]_net_1\, B => 
        \CONFIG_reg_14[3]_net_1\, C => un789_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(14), Y => 
        \edge_pos_147_iv_i_0[14]\);
    
    \edge_both_RNO[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[29]\, B => \CONFIG_reg_29[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(29), Y => 
        \edge_neg_297[29]\);
    
    \edge_neg_RNO[8]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[8]_net_1\, B => N_65, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        N_37_0);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_18\ : CFG3
      generic map(INIT => x"80")

      port map(A => un9_psel, B => m18_0, C => CONFIG_rega4, Y
         => un127_psel);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_5\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un156_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_5);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_8\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un242_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_8);
    
    edge_both_2_sqmuxa_440_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_14[3]_net_1\, D => un827_fixed_config, Y => 
        edge_both_2_sqmuxa_440_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_25\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un735_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_25);
    
    \GEN_BITS.11.APB_32.edge_neg_117_iv_i_RNO[11]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[11]_net_1\, B => 
        \CONFIG_reg_11[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(11), Y => N_183);
    
    \CONFIG_reg_17[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un503_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_17[6]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega25_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega25_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega23_2\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega23_2);
    
    g0_1_0 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \g0_1\);
    
    \edge_neg[17]\ : SLE
      port map(D => \edge_neg_177_iv_i_0[17]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_425_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[17]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_21\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un619_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_21);
    
    g0_1_0_a3_1 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \g0_1_0_a3_1\);
    
    \CONFIG_reg_2[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un69_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_2[3]_net_1\);
    
    \CONFIG_reg_14[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un416_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_14[5]_net_1\);
    
    \GPOUT_reg_RNII0ML5[6]\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \un30_psel\, B => m28_am_1, C => 
        \GPOUT_reg[6]_net_1\, Y => \GPOUT_reg_RNII0ML5[6]_net_1\);
    
    \CONFIG_reg_5[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un156_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_5[6]_net_1\);
    
    \GEN_BITS.14.APB_32.un827_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[14]_net_1\, B => \gpin3[14]_net_1\, Y
         => un827_fixed_config);
    
    \CONFIG_reg_18[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un532_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_18[5]_net_1\);
    
    \GEN_BITS.7.APB_32.edge_neg_77_iv_i_RNO[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[7]_net_1\, B => 
        \CONFIG_reg_7[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(7), Y => N_6192);
    
    \INTR_reg[28]\ : SLE
      port map(D => \INTR_reg_287[28]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[28]_net_1\);
    
    \CONFIG_reg_17[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un503_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_17[3]_net_1\);
    
    \GEN_BITS.1.REG_GPOUT.GPIO_OUT_i_3[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG_reg_1[0]_net_1\, B => 
        \GPOUT_reg[1]_net_1\, Y => GPIO_OUT_c(1));
    
    \edge_both_RNO[25]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[25]\, B => \CONFIG_reg_25[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(25), Y => 
        \edge_neg_257[25]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \INTR_reg_RNO_1[19]\ : CFG4
      generic map(INIT => x"8022")

      port map(A => \CONFIG_reg_19[3]_net_1\, B => m58_1_ns_1, C
         => \edge_both[19]_net_1\, D => \CONFIG_reg_19[7]_net_1\, 
        Y => N_59_0);
    
    \INTR_reg_RNO_0[7]\ : CFG4
      generic map(INIT => x"75FD")

      port map(A => \CONFIG_reg_7[3]_net_1\, B => 
        \CONFIG_reg_7[7]_net_1\, C => \INTR_reg_RNO_1[7]_net_1\, 
        D => m81_ns_1, Y => N_6158);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega21_0\ : CFG3
      generic map(INIT => x"20")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega21_0);
    
    \CONFIG_reg_15[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un445_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_15[5]_net_1\);
    
    \gpin1[4]\ : SLE
      port map(D => GPIO_IN_c(4), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[4]_net_1\);
    
    \edge_pos[17]\ : SLE
      port map(D => \edge_pos_177_iv_i_0[17]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_390_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[17]_net_1\);
    
    \INTR_reg_RNO[16]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[16]_net_1\, B => N_138_0, C => 
        CoreAPB3_0_APBmslave0_PWDATA(16), D => N_65, Y => 
        \INTR_reg_167[16]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_0_RNIRKRN1\ : CFG4
      generic map(INIT => x"C480")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        g0_6_a3_0, C => CONFIG_regro_4, D => CONFIG_regro_0, Y
         => g0_6_a3_2);
    
    \CONFIG_reg_11[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un329_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_11[3]_net_1\);
    
    \CONFIG_reg_0[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un11_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_0[7]_net_1\);
    
    m27_0 : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \m22_0_2\, D => 
        un1_psel_280_2, Y => un15_fixed_config);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_31_RNI1O5U1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega12_1, B => \CONFIG_rega23_1\, C
         => CONFIG_regro_31, D => CoreAPB3_0_APBmslave0_PADDR(6), 
        Y => CONFIG_regria_31);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_4\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega30_1, B => CONFIG_rega8_0, C => 
        m18_0, D => un9_psel, Y => un416_psel);
    
    \GEN_BITS.8.APB_32.edge_pos_87_iv_i[8]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[8]_net_1\, B => N_25_0, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        \edge_pos_87_iv_i_0[8]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_11_RNIVL5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega11_2, B => \CONFIG_rega23_1\, C
         => CONFIG_regro_11, D => CoreAPB3_0_APBmslave0_PADDR(6), 
        Y => CONFIG_regria_11);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega28_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega28_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega24_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => CONFIG_rega24_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_5_RNI3IN01\ : CFG3
      generic map(INIT => x"80")

      port map(A => CONFIG_regro_5, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => CONFIG_regria_5_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_10_RNIUL5U1\ : CFG4
      generic map(INIT => x"0400")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => g0_5_1, Y => 
        CONFIG_regria_10);
    
    \gpin3[9]\ : SLE
      port map(D => \gpin2[9]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[9]_net_1\);
    
    \edge_both_RNO_0[28]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_28[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_394_i_0);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNI8NPJ22\ : 
        CFG4
      generic map(INIT => x"3373")

      port map(A => \CONFIG_regror_29\, B => m57_ns_1, C => 
        m62_s_net_1, D => \CONFIG_regror_28\, Y => N_58);
    
    \edge_both_RNO[30]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[30]\, B => \CONFIG_reg_30[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(30), Y => 
        \edge_neg_307[30]\);
    
    \GEN_BITS.6.APB_32.edge_neg_67_iv_i_RNO[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[6]_net_1\, B => 
        \CONFIG_reg_6[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(6), Y => N_69_0);
    
    \CONFIG_reg_10_RNI10048[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_10[1]_net_1\, B => 
        \gpin3[10]_net_1\, C => \un3_prdata_o\, D => m357_ns_1, Y
         => N_358);
    
    \GEN_BITS.18.APB_32.edge_pos_187_iv_i[18]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[18]_net_1\, B => N_104_0, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        \edge_pos_187_iv_i_0[18]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega16_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega16_0);
    
    edge_neg_2_sqmuxa_409_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[6]_net_1\, B => N_65, C => 
        \gpin3[6]_net_1\, D => \CONFIG_reg_6[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_409_i_0);
    
    \CONFIG_reg_31[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un909_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_31[0]_net_1\);
    
    \CONFIG_reg_24[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un706_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_24[7]_net_1\);
    
    \GPOUT_reg[18]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(18), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[18]_net_1\);
    
    \GPOUT_reg[12]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(12), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[12]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_19_RNI7M5U1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega0_2, B => \CONFIG_rega23_1\, C => 
        CONFIG_regro_19, D => CoreAPB3_0_APBmslave0_PADDR(6), Y
         => CONFIG_regria_19);
    
    \CONFIG_reg_0[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un11_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_0[5]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega7\ : CFG4
      generic map(INIT => x"0200")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => \CONFIG_rega23_1\, Y
         => CONFIG_rega7);
    
    \GEN_BITS.11.APB_32.edge_both_117_iv_i[11]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[11]_net_1\, B => 
        \CONFIG_reg_11[3]_net_1\, C => un659_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(11), Y => 
        \edge_both_117_iv_i_0[11]\);
    
    \CONFIG_reg_16[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un474_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_16[5]_net_1\);
    
    \CONFIG_reg_16[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un474_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_16[1]_net_1\);
    
    \GEN_BITS.13.APB_32.edge_both_137_iv_i[13]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[13]_net_1\, B => N_201, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        \edge_both_137_iv_i_0[13]\);
    
    \CONFIG_reg_15[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un445_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_15[7]_net_1\);
    
    \GEN_BITS.23.APB_32.INTR_reg_237_ns[23]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(23), B => N_65, 
        C => \INTR_reg[23]_net_1\, D => \INTR_reg_237_ns_1[23]\, 
        Y => \INTR_reg_237[23]\);
    
    \edge_both_RNO[2]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[2]\, B => \CONFIG_reg_2[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(2), Y => 
        \edge_neg_27[2]\);
    
    \GPOUT_reg[28]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(28), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_28);
    
    \edge_both_RNO[31]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[31]\, B => \CONFIG_reg_31[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(31), Y => 
        \edge_neg_317[31]\);
    
    \edge_both_RNO[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_pos[26]\, B => \CONFIG_reg_26[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(26), Y => 
        \edge_neg_267[26]\);
    
    \INTR_reg[24]\ : SLE
      port map(D => \INTR_reg_247[24]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[24]_net_1\);
    
    \GPOUT_reg[22]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(22), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_22);
    
    \GEN_BITS.5.APB_32.edge_both_57_iv_i[5]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[5]_net_1\, B => N_6152, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        \edge_both_57_iv_i_0[5]\);
    
    g0_2_1 : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \g0_2_1\);
    
    g0_1_0_a3 : CFG4
      generic map(INIT => x"0010")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \g0_1_0_a3_1\, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega0);
    
    \edge_both_RNO_0[9]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[9]_net_1\, B => N_65, C => 
        \gpin3[9]_net_1\, D => \CONFIG_reg_9[3]_net_1\, Y => 
        \edge_both_RNO_0[9]_net_1\);
    
    \CONFIG_reg_19[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un561_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_19[7]_net_1\);
    
    \GEN_BITS.11.APB_32.edge_neg_117_iv_i[11]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[11]_net_1\, B => N_183, C => 
        \gpin3[11]_net_1\, D => \CONFIG_reg_11[3]_net_1\, Y => 
        \edge_neg_117_iv_i_0[11]\);
    
    \CONFIG_reg_16[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un474_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_16[7]_net_1\);
    
    \CONFIG_reg_12[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un358_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_12[3]_net_1\);
    
    \INTR_reg_RNO_0[14]\ : CFG4
      generic map(INIT => x"C480")

      port map(A => \CONFIG_reg_14[6]_net_1\, B => 
        \CONFIG_reg_14[3]_net_1\, C => \INTR_reg_RNO_1[14]_net_1\, 
        D => \INTR_reg_RNO_2[14]_net_1\, Y => N_6250);
    
    \CONFIG_reg_2[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un69_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_2[7]_net_1\);
    
    \CONFIG_reg_10[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un300_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_10[6]_net_1\);
    
    edge_pos_2_sqmuxa_375_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_4[3]_net_1\, D => un229_fixed_config, Y => 
        edge_pos_2_sqmuxa_375_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_28_RNI7N5U1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CONFIG_rega12_1, B => CONFIG_rega26_2, C => 
        CONFIG_regro_28, D => CoreAPB3_0_APBmslave0_PADDR(3), Y
         => CONFIG_regria_28);
    
    \CONFIG_reg_4[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un127_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_4[7]_net_1\);
    
    \gpin3[17]\ : SLE
      port map(D => \gpin2[17]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[17]_net_1\);
    
    \GPOUT_reg_RNIREG25[14]\ : CFG4
      generic map(INIT => x"15BF")

      port map(A => \N_6186\, B => \un30_psel\, C => 
        \GPOUT_reg[14]_net_1\, D => \INTR_reg[14]_net_1\, Y => 
        m318_ns_1);
    
    \CONFIG_reg_12[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un358_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_12[1]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNO\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => un9_psel, B => m18_0, Y => CONFIG_reg_0_0_we);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_10\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un300_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_10);
    
    \CONFIG_reg_10[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un300_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_10[7]_net_1\);
    
    \gpin1[14]\ : SLE
      port map(D => GPIO_IN_c(14), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[14]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_29\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un851_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_29);
    
    \CONFIG_reg_30[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un880_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_30[5]_net_1\);
    
    \CONFIG_reg_17[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un503_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_17[7]_net_1\);
    
    \edge_pos[13]\ : SLE
      port map(D => \edge_pos_137_iv_i_0[13]\, CLK => FAB_CCC_GL0, 
        EN => N_216, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_pos[13]_net_1\);
    
    \CONFIG_reg_4_RNII8VS2[1]\ : CFG4
      generic map(INIT => x"35F5")

      port map(A => \INTR_reg[4]_net_1\, B => 
        \CONFIG_reg_4[1]_net_1\, C => \un3_prdata_o\, D => 
        \gpin3[4]_net_1\, Y => m41_am_1);
    
    g0_11 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => g0_1_2);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIIPJD8\ : 
        CFG4
      generic map(INIT => x"4073")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        m62_s_net_1, C => \CONFIG_regrx[6]\, D => 
        \GPOUT_reg_RNII0ML5[6]_net_1\, Y => N_122_i_1);
    
    \GEN_BITS.4.APB_32.edge_pos_47_iv_i[4]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_pos[4]_net_1\, B => 
        \CONFIG_reg_4[3]_net_1\, C => un229_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(4), Y => 
        \edge_pos_47_iv_i_0[4]\);
    
    \GEN_BITS.17.APB_32.edge_neg_177_iv_i[17]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_neg[17]_net_1\, B => 
        \CONFIG_reg_17[3]_net_1\, C => un977_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(17), Y => 
        \edge_neg_177_iv_i_0[17]\);
    
    \GEN_BITS.23.APB_32.INTR_reg_237_ns_1_1[23]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_23[5]_net_1\, B => \edge_neg[23]\, 
        C => \CONFIG_reg_23[7]_net_1\, D => 
        \CONFIG_reg_23[6]_net_1\, Y => \INTR_reg_237_ns_1_1[23]\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNI6LPJ22\ : 
        CFG4
      generic map(INIT => x"3373")

      port map(A => \CONFIG_regror_29\, B => m62_ns_1, C => 
        m62_s_net_1, D => \CONFIG_regror_28\, Y => N_63);
    
    \edge_neg_RNO[18]\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[18]_net_1\, B => N_65, C => 
        \gpin3[18]_net_1\, D => \CONFIG_reg_18[3]_net_1\, Y => 
        N_113_0);
    
    \edge_both_RNO_0[12]\ : CFG4
      generic map(INIT => x"7BFF")

      port map(A => \gpin2[12]_net_1\, B => N_65, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        \edge_both_RNO_0[12]_net_1\);
    
    \GEN_BITS.25.APB_32.INTR_reg_257_ns_1[25]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_257_ns_1_1[25]\, B => 
        \CONFIG_reg_25[3]_net_1\, Y => \INTR_reg_257_ns_1[25]\);
    
    \GEN_BITS.17.APB_32.un977_fixed_config\ : CFG2
      generic map(INIT => x"4")

      port map(A => \gpin2[17]_net_1\, B => \gpin3[17]_net_1\, Y
         => un977_fixed_config);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_11_RNIABEP8\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => CONFIG_regria_10, B => CONFIG_regria_26, C
         => CONFIG_regria_11, D => CONFIG_regror_0, Y => 
        CONFIG_regror_22);
    
    \GEN_BITS.30.APB_32.INTR_reg_307_ns_1[30]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_307_ns_1_1[30]\, B => 
        \CONFIG_reg_30[3]_net_1\, Y => \INTR_reg_307_ns_1[30]\);
    
    \CONFIG_reg_25[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un735_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_25[3]_net_1\);
    
    \edge_pos[8]\ : SLE
      port map(D => \edge_pos_87_iv_i_0[8]\, CLK => FAB_CCC_GL0, 
        EN => N_36_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \edge_pos[8]_net_1\);
    
    \CONFIG_reg_6[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un185_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_6[7]_net_1\);
    
    \CONFIG_reg_12[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un358_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_12[5]_net_1\);
    
    \gpin3[15]\ : SLE
      port map(D => \gpin2[15]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[15]_net_1\);
    
    \gpin2[10]\ : SLE
      port map(D => \gpin1[10]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[10]_net_1\);
    
    \edge_both[9]\ : SLE
      port map(D => i21_mux, CLK => FAB_CCC_GL0, EN => 
        \edge_both_RNO_0[9]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[9]_net_1\);
    
    \GEN_BITS.26.APB_32.INTR_reg_267_ns_1[26]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \INTR_reg_267_ns_1_1[26]\, B => 
        \CONFIG_reg_26[3]_net_1\, Y => \INTR_reg_267_ns_1[26]\);
    
    \CONFIG_reg_9[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un271_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_9[3]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_1_RNI7SRE1\ : CFG4
      generic map(INIT => x"3FF5")

      port map(A => CONFIG_regro_1, B => CONFIG_regro_13, C => 
        CoreAPB3_0_APBmslave0_PADDR(5), D => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => g0_0_1_1);
    
    \CONFIG_reg_17[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un503_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_17[5]_net_1\);
    
    \CONFIG_reg_15[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un445_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_15[6]_net_1\);
    
    \CONFIG_reg_22[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un648_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_22[6]_net_1\);
    
    \GEN_BITS.16.APB_32.un939_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[16]_net_1\, B => \gpin3[16]_net_1\, Y
         => un939_fixed_config);
    
    \CONFIG_reg_24[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un706_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_24[6]_net_1\);
    
    \CONFIG_reg_16_RNIP4JQ7[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_16[1]_net_1\, B => 
        \gpin3[16]_net_1\, C => \un3_prdata_o\, D => m327_ns_1, Y
         => N_328);
    
    \GEN_BITS.14.APB_32.edge_both_147_iv_i[14]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[14]_net_1\, B => 
        \CONFIG_reg_14[3]_net_1\, C => un827_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(14), Y => 
        \edge_both_147_iv_i_0[14]\);
    
    \CONFIG_reg_20[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un590_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_20[3]_net_1\);
    
    \INTR_reg_RNITM6H2[29]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[29]_net_1\, Y => INTR_reg_m_7);
    
    \CONFIG_reg_29[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un851_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_29[5]_net_1\);
    
    \GPOUT_reg[14]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(14), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \GPOUT_reg[14]_net_1\);
    
    \gpin2[18]\ : SLE
      port map(D => \gpin1[18]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin2[18]_net_1\);
    
    edge_neg_2_sqmuxa_408_i : CFG4
      generic map(INIT => x"73FF")

      port map(A => \gpin2[7]_net_1\, B => N_65, C => 
        \gpin3[7]_net_1\, D => \CONFIG_reg_7[3]_net_1\, Y => 
        edge_neg_2_sqmuxa_408_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regwre_23\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CONFIG_rega23_2, C => \CONFIG_rega23_1\, D => 
        un11_psel_1_0, Y => un677_psel);
    
    \GEN_BITS.8.APB_32.edge_both_87_iv_i[8]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[8]_net_1\, B => N_6244, C => 
        \gpin3[8]_net_1\, D => \CONFIG_reg_8[3]_net_1\, Y => 
        \edge_both_87_iv_i_0[8]\);
    
    \edge_both_RNO_1[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_both[10]_net_1\, B => 
        \CONFIG_reg_10[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(10), Y => N_292);
    
    \edge_both[10]\ : SLE
      port map(D => i15_mux, CLK => FAB_CCC_GL0, EN => 
        \edge_both_RNO_0[10]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_both[10]_net_1\);
    
    \INTR_reg_RNO[0]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[0]_net_1\, B => N_6170, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), D => N_65, Y => 
        N_6172_i_0);
    
    \GPOUT_reg[24]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(24), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_24);
    
    \CONFIG_reg_23[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un677_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_23[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega18\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => CONFIG_rega18_1, Y
         => CONFIG_rega18);
    
    \CONFIG_reg_10[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un300_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_10[1]_net_1\);
    
    \INTR_reg_RNO_0[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_6177, B => \CONFIG_reg_1[3]_net_1\, Y => 
        \intr_3[1]\);
    
    \CONFIG_reg_12[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un358_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_12[7]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIAPPJ22\ : 
        CFG4
      generic map(INIT => x"3373")

      port map(A => \CONFIG_regror_29\, B => m52_ns_1, C => 
        m62_s_net_1, D => \CONFIG_regror_28\, Y => N_53);
    
    \edge_pos_RNO[13]\ : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[13]_net_1\, B => N_65, C => 
        \gpin3[13]_net_1\, D => \CONFIG_reg_13[3]_net_1\, Y => 
        N_216);
    
    \edge_both_RNO_0[25]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_25[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_382_i_0);
    
    \edge_both[31]\ : SLE
      port map(D => \edge_neg_317[31]\, CLK => FAB_CCC_GL0, EN
         => edge_neg_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[31]\);
    
    \INTR_reg[8]\ : SLE
      port map(D => \INTR_reg_87[8]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[8]_net_1\);
    
    \INTR_reg_RNIRK6H2[27]\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => \N_6186\, 
        C => \INTR_reg[27]_net_1\, Y => N_441);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega12_1, B => CONFIG_rega0_0, C => 
        un9_psel, D => m18_0, Y => un358_psel);
    
    \edge_pos[4]\ : SLE
      port map(D => \edge_pos_47_iv_i_0[4]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_375_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[4]_net_1\);
    
    \INTR_reg_RNO_3[18]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_18[6]_net_1\, B => 
        \edge_pos[18]_net_1\, C => \gpin3[18]_net_1\, D => 
        \CONFIG_reg_18[7]_net_1\, Y => m93_0_ns_1);
    
    \GEN_BITS.24.APB_32.INTR_reg_247_ns[24]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(24), B => N_65, 
        C => \INTR_reg[24]_net_1\, D => \INTR_reg_247_ns_1[24]\, 
        Y => \INTR_reg_247[24]\);
    
    \edge_both_RNO_0[27]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_27[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_395_i_0);
    
    \CONFIG_reg_8[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un242_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_8[1]_net_1\);
    
    \gpin1[16]\ : SLE
      port map(D => GPIO_IN_c(16), CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin1[16]_net_1\);
    
    \edge_both_RNO_0[21]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_21[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_400_i_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_3_RNIT23O7\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => CONFIG_regria_27, B => CONFIG_regria_16, C
         => CONFIG_regria_3, D => CONFIG_regria_15, Y => 
        CONFIG_regror_18);
    
    \CONFIG_reg_28[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un822_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_28[3]_net_1\);
    
    \INTR_reg_RNO[6]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[6]_net_1\, B => m50_0_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(6), D => N_65, Y => 
        \INTR_reg_67[6]\);
    
    \INTR_reg[27]\ : SLE
      port map(D => \INTR_reg_277[27]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[27]_net_1\);
    
    \INTR_reg_RNO_3[6]\ : CFG4
      generic map(INIT => x"5527")

      port map(A => \CONFIG_reg_6[6]_net_1\, B => 
        \edge_pos[6]_net_1\, C => \gpin3[6]_net_1\, D => 
        \CONFIG_reg_6[7]_net_1\, Y => m44_1_ns_1);
    
    \INTR_reg[25]\ : SLE
      port map(D => \INTR_reg_257[25]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[25]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_10_RNIF8B11\ : CFG3
      generic map(INIT => x"20")

      port map(A => CONFIG_regro_10, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => g0_5_1);
    
    \edge_both_RNO[3]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[3]\, B => \CONFIG_reg_3[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \edge_neg_37[3]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega17\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), D => CONFIG_rega17_1, Y
         => CONFIG_rega17);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega11_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => CONFIG_rega11_2);
    
    \CONFIG_reg_12_RNIERPV7[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_12[1]_net_1\, B => 
        \gpin3[12]_net_1\, C => \un3_prdata_o\, D => m309_ns_1, Y
         => N_310);
    
    \CONFIG_reg_29[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un851_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_29[6]_net_1\);
    
    \INTR_reg_RNO_1[7]\ : CFG4
      generic map(INIT => x"EB41")

      port map(A => \CONFIG_reg_7[6]_net_1\, B => 
        \CONFIG_reg_7[5]_net_1\, C => \gpin3[7]_net_1\, D => 
        N_6193, Y => \INTR_reg_RNO_1[7]_net_1\);
    
    \INTR_reg_RNO_1[2]\ : CFG4
      generic map(INIT => x"0C4A")

      port map(A => \CONFIG_reg_2[5]_net_1\, B => \edge_neg[2]\, 
        C => \CONFIG_reg_2[7]_net_1\, D => 
        \CONFIG_reg_2[6]_net_1\, Y => m67_0_ns_1_0);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega3_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega3_0);
    
    INTR_reg_0_sqmuxa_0_o2 : CFG3
      generic map(INIT => x"DF")

      port map(A => un9_psel, B => CoreAPB3_0_APBmslave0_PADDR(4), 
        C => \N_6186\, Y => N_65);
    
    g0_14 : CFG3
      generic map(INIT => x"08")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega9_0);
    
    \GPOUT_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => N_51_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => GPOUT_reg_3);
    
    \edge_pos[5]\ : SLE
      port map(D => \edge_pos_57_iv_i_0[5]\, CLK => FAB_CCC_GL0, 
        EN => edge_pos_2_sqmuxa_389_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_pos[5]_net_1\);
    
    edge_neg_2_sqmuxa_425_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_17[3]_net_1\, D => un977_fixed_config, Y => 
        edge_neg_2_sqmuxa_425_i_0);
    
    \INTR_reg_RNO_1[14]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => \edge_pos[14]_net_1\, B => 
        \edge_neg[14]_net_1\, C => \CONFIG_reg_14[7]_net_1\, D
         => \CONFIG_reg_14[5]_net_1\, Y => 
        \INTR_reg_RNO_1[14]_net_1\);
    
    \CONFIG_reg_8[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un242_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_8[5]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega16_2, B => CONFIG_rega8_0, C => 
        m18_0, D => un9_psel, Y => un242_psel);
    
    \CONFIG_reg_11[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un329_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_11[5]_net_1\);
    
    \INTR_reg_RNO[9]\ : CFG4
      generic map(INIT => x"330A")

      port map(A => \INTR_reg[9]_net_1\, B => m244_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(9), D => N_65, Y => 
        \INTR_reg_97[9]\);
    
    \GEN_BITS.31.APB_32.INTR_reg_317_ns[31]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(31), B => N_65, 
        C => \INTR_reg[31]_net_1\, D => \INTR_reg_317_ns_1[31]\, 
        Y => \INTR_reg_317[31]\);
    
    \INTR_reg_RNO_3[12]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => \edge_neg[12]_net_1\, B => 
        \edge_pos[12]_net_1\, C => \CONFIG_reg_12[6]_net_1\, D
         => \CONFIG_reg_12[5]_net_1\, Y => m269_ns_1);
    
    \edge_pos_RNO[10]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[10]_net_1\, B => N_282, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        N_44);
    
    \CONFIG_reg_11[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un329_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_11[7]_net_1\);
    
    \INTR_reg[5]\ : SLE
      port map(D => N_92_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \INTR_reg[5]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_31\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un909_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_31);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_6_RNIA8JUU\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => CONFIG_regror_29_1, B => CONFIG_regror_23, C
         => CONFIG_regror_22, D => CONFIG_regror_11, Y => 
        \CONFIG_regror_29\);
    
    \edge_both[24]\ : SLE
      port map(D => \edge_neg_247[24]\, CLK => FAB_CCC_GL0, EN
         => edge_pos_2_sqmuxa_397_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[24]\);
    
    \GEN_BITS.11.APB_32.un659_fixed_config\ : CFG2
      generic map(INIT => x"6")

      port map(A => \gpin2[11]_net_1\, B => \gpin3[11]_net_1\, Y
         => un659_fixed_config);
    
    \CONFIG_reg_18_RNI60D68[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_18[1]_net_1\, B => 
        \gpin3[18]_net_1\, C => \un3_prdata_o\, D => m337_ns_1, Y
         => N_338);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_17_RNI3JFF1\ : CFG4
      generic map(INIT => x"0CA0")

      port map(A => CONFIG_regro_18, B => CONFIG_regro_17, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        CONFIG_regrff_17_RNI3JFF1);
    
    \GEN_BITS.4.APB_32.edge_both_47_iv_i[4]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[4]_net_1\, B => 
        \CONFIG_reg_4[3]_net_1\, C => un267_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(4), Y => 
        \edge_both_47_iv_i_0[4]\);
    
    \gpin3[19]\ : SLE
      port map(D => \gpin2[19]_net_1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \gpin3[19]_net_1\);
    
    
        \GEN_BITS.0.REG_GEN.CONFIG_reg_GEN_BITS.0.REG_GEN.CONFIG_reg_0_0_RNIOTH78\ : 
        CFG4
      generic map(INIT => x"2075")

      port map(A => m62_s_net_1, B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => \CONFIG_regrx[1]\, D
         => \GPOUT_reg_RNIO4KF5[1]_net_1\, Y => m57_ns_1);
    
    edge_pos_2_sqmuxa_389_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[5]_net_1\, B => N_65, C => 
        \gpin3[5]_net_1\, D => \CONFIG_reg_5[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_389_i_0);
    
    \CONFIG_reg_4[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un127_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_4[5]_net_1\);
    
    edge_pos_2_sqmuxa_379_i : CFG4
      generic map(INIT => x"FF8F")

      port map(A => un15_fixed_config, B => un9_psel, C => 
        \CONFIG_reg_14[3]_net_1\, D => un789_fixed_config, Y => 
        edge_pos_2_sqmuxa_379_i_0);
    
    \CONFIG_reg_13[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un387_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_13[6]_net_1\);
    
    \CONFIG_reg_6[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un185_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_6[5]_net_1\);
    
    \INTR_reg[23]\ : SLE
      port map(D => \INTR_reg_237[23]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[23]_net_1\);
    
    \GEN_BITS.22.APB_32.INTR_reg_227_ns[22]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(22), B => N_65, 
        C => \INTR_reg[22]_net_1\, D => \INTR_reg_227_ns_1[22]\, 
        Y => \INTR_reg_227[22]\);
    
    \INTR_reg_RNO_2[18]\ : CFG4
      generic map(INIT => x"3FBB")

      port map(A => \gpin3[18]_net_1\, B => 
        \CONFIG_reg_18[3]_net_1\, C => \edge_neg[18]_net_1\, D
         => \CONFIG_reg_18[6]_net_1\, Y => N_97_0);
    
    \CONFIG_reg_1[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un41_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_1[0]_net_1\);
    
    \CONFIG_reg_19[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un561_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_19[1]_net_1\);
    
    g0_2 : CFG4
      generic map(INIT => x"0080")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \g0_2_1\, D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => CONFIG_rega13);
    
    \CONFIG_reg_5[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un156_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_5[7]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_12\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega30_2, B => CONFIG_rega24_0, C => 
        un9_psel, D => m18_0, Y => un706_psel);
    
    \GEN_BITS.6.APB_32.edge_pos_67_iv_i[6]\ : CFG4
      generic map(INIT => x"CEC4")

      port map(A => \gpin2[6]_net_1\, B => N_75_0, C => 
        \gpin3[6]_net_1\, D => \CONFIG_reg_6[3]_net_1\, Y => 
        \edge_pos_67_iv_i_0[6]\);
    
    \CONFIG_reg_5[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un156_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_5[3]_net_1\);
    
    edge_pos_2_sqmuxa_402_i : CFG4
      generic map(INIT => x"3BFF")

      port map(A => \gpin2[19]_net_1\, B => N_65, C => 
        \gpin3[19]_net_1\, D => \CONFIG_reg_19[3]_net_1\, Y => 
        edge_pos_2_sqmuxa_402_i_0);
    
    \edge_neg_RNO[12]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[12]_net_1\, B => N_279, C => 
        \gpin3[12]_net_1\, D => \CONFIG_reg_12[3]_net_1\, Y => 
        N_46);
    
    \GPOUT_reg_RNI864C5[18]\ : CFG4
      generic map(INIT => x"353F")

      port map(A => \GPOUT_reg[18]_net_1\, B => 
        \INTR_reg[18]_net_1\, C => un15_fixed_config, D => 
        \un30_psel\, Y => m337_ns_1);
    
    \INTR_reg_RNO[13]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[13]_net_1\, B => m167_ns_1, C => 
        CoreAPB3_0_APBmslave0_PWDATA(13), D => N_65, Y => 
        \INTR_reg_137[13]\);
    
    \edge_both_RNO[10]\ : CFG4
      generic map(INIT => x"DE84")

      port map(A => \gpin2[10]_net_1\, B => N_292, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        i15_mux);
    
    \CONFIG_reg_7[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un214_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_7[3]_net_1\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_regrff_20\ : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        un590_psel, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CONFIG_regro_20);
    
    \edge_both_RNO_0[2]\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \CONFIG_reg_2[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => \N_6186\, D => 
        un9_psel, Y => edge_pos_2_sqmuxa_378_i_0);
    
    \INTR_reg_RNO_2[12]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \edge_both[12]_net_1\, B => 
        \CONFIG_reg_12[5]_net_1\, C => \CONFIG_reg_12[6]_net_1\, 
        D => \CONFIG_reg_12[3]_net_1\, Y => N_434_mux);
    
    \INTR_reg_RNO[5]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => \INTR_reg[5]_net_1\, B => N_90, C => 
        CoreAPB3_0_APBmslave0_PWDATA(5), D => N_65, Y => N_92_i_0);
    
    \INTR_reg[11]\ : SLE
      port map(D => \INTR_reg_117[11]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INTR_reg[11]_net_1\);
    
    \edge_neg[15]\ : SLE
      port map(D => \edge_neg_157_iv_i_0[15]\, CLK => FAB_CCC_GL0, 
        EN => edge_neg_2_sqmuxa_427_i_0, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \edge_neg[15]_net_1\);
    
    \GEN_BITS.0.REG_GEN.un9_psel_RNIB00P2_2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CONFIG_rega21_1, B => CONFIG_rega5_0, C => 
        m18_0, D => un9_psel, Y => un156_psel);
    
    \CONFIG_reg_14_RNIHOCO7[1]\ : CFG4
      generic map(INIT => x"7F70")

      port map(A => \CONFIG_reg_14[1]_net_1\, B => 
        \gpin3[14]_net_1\, C => \un3_prdata_o\, D => m318_ns_1, Y
         => N_319);
    
    \GEN_BITS.6.APB_32.edge_neg_67_iv_i[6]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[6]_net_1\, B => N_69_0, C => 
        \gpin3[6]_net_1\, D => \CONFIG_reg_6[3]_net_1\, Y => 
        \edge_neg_67_iv_i_0[6]\);
    
    \GEN_BITS.16.APB_32.edge_both_167_iv_i[16]\ : CFG4
      generic map(INIT => x"C0C8")

      port map(A => \edge_both[16]_net_1\, B => 
        \CONFIG_reg_16[3]_net_1\, C => un939_fixed_config, D => 
        CoreAPB3_0_APBmslave0_PWDATA(16), Y => 
        \edge_both_167_iv_i_0[16]\);
    
    \CONFIG_reg_11[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un329_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_11[6]_net_1\);
    
    \GEN_BITS.16.APB_32.un901_fixed_config\ : CFG2
      generic map(INIT => x"2")

      port map(A => \gpin2[16]_net_1\, B => \gpin3[16]_net_1\, Y
         => un901_fixed_config);
    
    g0_5_0_a3_1 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \g0_5_0_a3_1\);
    
    \edge_neg_RNO[10]\ : CFG4
      generic map(INIT => x"DC8C")

      port map(A => \gpin2[10]_net_1\, B => N_276, C => 
        \gpin3[10]_net_1\, D => \CONFIG_reg_10[3]_net_1\, Y => 
        N_48);
    
    \edge_both_RNO[23]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \edge_neg[23]\, B => \CONFIG_reg_23[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PWDATA(23), Y => 
        \edge_neg_237[23]\);
    
    \GEN_BITS.0.REG_GEN.CONFIG_rega30_2\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => CONFIG_rega30_2);
    
    \CONFIG_reg_3[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un98_psel, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \CONFIG_reg_3[7]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6 is

    port( COREI2C_0_0_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0);
          seradr0apb                                 : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          CONFIG_rega20_2                            : out   std_logic;
          bclke                                      : in    std_logic;
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_0_SDA_IO_Y                 : in    std_logic;
          un105_ens1_3                               : out   std_logic;
          BIBUF_COREI2C_0_0_SCL_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          un3_penable_1                              : out   std_logic;
          un5_penable_0                              : out   std_logic;
          un105_ens1_0                               : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_138                                      : in    std_logic;
          un5_penable_2                              : in    std_logic
        );

end COREI2CREAL_6;

architecture DEF_ARCH of COREI2CREAL_6 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_0_SDAO[0]\, \COREI2C_0_0_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_0_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        \un1_serdat_2_sqmuxa\, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, fsmsta_8_5_555, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, fsmsta_8_28_307, \ack\, ack_7, N_1449, 
        SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, bsd7_tmp_6, \bsd7\, 
        bsd7_9_iv_i_0, \adrcomp\, N_2176, \adrcomp_2_sqmuxa_i_0\, 
        \PCLKint\, PCLKint_3, un1_pclkint4_i_0, \ack_bit\, 
        \ack_bit_1_sqmuxa\, \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        \un1_rtn_4\, \un1_rtn_3\, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, PCLK_count2_ov_6_1, 
        \PCLK_count1_1_sqmuxa_1\, CO1, N_126, N_2181, 
        un133_framesync, N_80, N_2199, N_157, un70_fsmsta, CO0, 
        N_1586_1, N_1656, \fsmsta_cnst[0]\, N_2188, N_2177, 
        N_2179, N_162, \adrcomp_2_sqmuxa_i_o2_1_3\, un57_fsmsta_0, 
        un57_fsmsta_1_0, un57_fsmsta, N_2173_i_1, un1_fsmmod, 
        N_133, N_36_i_1, un136_framesync, N_2196, N_2186, 
        \fsmsta_8_1[24]\, N_172, fsmsta_8_3_601_0_1, N_1717, 
        fsmsta_8_3_601_0, N_1652, fsmsta_8_9_509_0_1, 
        fsmsta_8_9_509_0, \un1_pclk_count1_ov_1_1\, 
        \un1_pclk_count1_ov_1\, \PCLK_count1_1_sqmuxa_1_0_1\, 
        \PCLK_count1_1_sqmuxa_1_0\, CO1_0, \PRDATA_3_1_1[7]\, 
        \PRDATA_3_1_1[3]\, \PRDATA_3_1_1[6]\, \PRDATA_3_1_1[4]\, 
        \PRDATA_3_1_1[5]\, \fsmsta_8_ns_1[29]\, 
        \fsmsta_8_ns_1[28]\, \fsmsta_8_ns_1[18]\, un13_adrcompen, 
        \fsmsta_8_ns_1[16]\, bsd7_tmp_6_am, bsd7_tmp_6_ns_1, 
        un92_fsmsta, un105_ens1, N_161_2, fsmsta_8_5_555_a3_2, 
        fsmsta_8_5_555_a3_0_2, PCLK_count2_ov_6_0_a2_1_0, 
        \fsmsta_nxt_9_m_0[26]\, \fsmsta_nxt_9_m_0[21]\, 
        \sersta_32_2[0]\, un111_fsmdet_0, \sersta_32_i_a2_5[3]\, 
        \PCLK_count1_ov_1_sqmuxa_0\, un139_ens1_0, 
        fsmsta_8_20_379_i_0_a3_3, \adrcomp_2_sqmuxa_i_o2_1_1\, 
        un135_ens1_7, N_26, N_127, N_23, N_2178, \un1_fsmsta_2_1\, 
        N_64, N_1035, N_67, N_1002_3, \un151_framesync\, 
        un26_adrcompen_6, \un105_ens1_3\, N_145_2, N_1196, N_1197, 
        N_1198, SDAO_int_7_0_275_1, \adrcomp_2_sqmuxa_i_a3_3\, 
        SDAO_int_7_0_275_a5_0, un141_ens1_2, 
        \SDAO_int_1_sqmuxa_3\, \adrcomp_2_sqmuxa_i_a2_1_2\, 
        \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_10_476_i_a6_1, 
        \sersta_32_5[1]\, \sersta_32_4[1]\, \sersta_32_3[0]\, 
        fsmsta_8_20_379_i_0_a3_4, fsmsta_8_20_379_i_0_a3_3_0, 
        \sersta_32_i_a2_7[4]\, \sersta_32_i_a2_6[4]\, 
        \sersta_32_6[2]\, \sersta_32_4[2]\, un135_ens1_4, 
        un135_ens1_3, fsmsta_nxt_1_sqmuxa_24_s4_1_0, 
        un25_fsmsta_1, \sersta_32_i_a2_8[3]\, 
        \sersta_32_i_a2_7[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, m7_3, 
        \PCLK_count1_0_sqmuxa_4_1\, un13_adrcompen_4, 
        \un3_penable_1\, un33_fsmsta, framesync_7_e2_1, N_1064, 
        \un105_ens1_0\, PCLK_count2_ov_6_0_a2_1_4_tz, N_1034, 
        N_2182, N_1049, N_68, N_1040, N_76, N_189, N_163_2, ANC2, 
        CO2, \un1_pclk_count1_ov\, CO1_1, N_95, un16_fsmmod, 
        \adrcomp_2_sqmuxa_i_a3_4\, \fsmmod_ns_i_0[2]_net_1\, 
        fsmsta_8_10_476_i_0, \SDAO_int_1_sqmuxa_4\, 
        \fsmsync_ns_i_0[6]_net_1\, \adrcomp_2_sqmuxa_i_a2_1_4\, 
        PCLK_count2_ov_6_0_a2_1_3, \fsmmod_ns_i_a4_1_1[2]_net_1\, 
        \sercon_8_2[4]\, \sersta_32_i_a2_9[4]\, \sersta_32_7[2]\, 
        un135_ens1_7_0, \sersta_32_i_a2_10[3]\, N_72_mux, N_104, 
        N_1002, N_2192, un19_framesync, un25_framesync, 
        fsmsta_nxt_1_sqmuxa_18_s5_1, un25_fsmsta, N_130, N_2193, 
        N_2171, un74_ens1, un8_nedetect, N_84, N_63, 
        \un1_fsmsta_6\, N_1622_2, \un1_pclk_count191\, un91_ens1, 
        N_124, N_120, fsmsta_8_28_307_a3_0_1, fsmsta_8_9_509_a4_0, 
        fsmsta_8_3_601_a4_0, \SDAO_int_1_sqmuxa_7\, 
        \adrcomp_2_sqmuxa_i_a2_1_5\, N_1007, un115_fsmdet, 
        \fsmsta_nxt_9_m[27]\, N_108, un135_ens1, 
        \PCLK_count1_0_sqmuxa_1\, \fsmsta_nxt_9_m[22]\, N_165, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, N_1046, N_193, N_1048, 
        N_1060, N_70, N_1624, \PCLK_count1_0_sqmuxa_2\, 
        \PCLK_count1_0_sqmuxa_3\, \fsmsta_8_i_0[25]\, 
        fsmsta_8_4_577_i_0, N_82, bsd7_tmp_i_m_2, 
        bsd7_tmp_6_sn_m6_1, fsmsta_8_20_379_i_0_o2_0, 
        \sercon_8_0_1[3]\, \sercon_8_0_0[3]\, 
        \fsmmod_ns_i_1[2]_net_1\, fsmsta_8_23_351_i_0_1, 
        \fsmsync_ns_0_0_1[0]_net_1\, 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\, N_1058, N_166, N_145, 
        N_1465, \fsmsync_ns_i_0_1_tz[3]_net_1\, N_1059_1, CO1_2, 
        N_86, \PWDATA_i_m_1[7]\, \PCLK_count1_1_sqmuxa_3\, 
        fsmsta_8_2_647_i_0_0, N_1486, N_1051, \framesync_7_m2[3]\, 
        framesync_7_e2, CO2_0, N_2187, \fsmsta_s12[21]\, 
        \serdat_0_sqmuxa\, un134_fsmsta, N_1466, \sercon_8[3]\, 
        \serdat_2_sqmuxa\, \un1_bsd7_1_sqmuxa[0]_net_1\, 
        \un1_serdat40\, bsd7_9_iv_1, \serdat_1_sqmuxa_1\, 
        \un1_counter_rst_3\, bsd7_9_iv_2, \un1_serdat_2_sqmuxa_1\
         : std_logic;

begin 

    COREI2C_0_0_INT(0) <= \COREI2C_0_0_INT[0]\;
    un105_ens1_3 <= \un105_ens1_3\;
    un3_penable_1 <= \un3_penable_1\;
    un105_ens1_0 <= \un105_ens1_0\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[21]\);
    
    \un1_bsd7_1_sqmuxa[0]\ : CFG3
      generic map(INIT => x"A1")

      port map(A => un105_ens1, B => \nedetect\, C => 
        \COREI2C_0_0_INT[0]\, Y => \un1_bsd7_1_sqmuxa[0]_net_1\);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    adrcomp_2_sqmuxa_i_0_0 : CFG4
      generic map(INIT => x"0015")

      port map(A => un16_fsmmod, B => N_2192, C => 
        \COREI2C_0_0_INT[0]\, D => N_1586_1, Y => N_2176);
    
    \fsmmod_RNIS2JA2[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_189, B => \fsmsta_cnst[0]\, Y => N_1622_2);
    
    \un2_framesync_1_1.CO2\ : CFG2
      generic map(INIT => x"8")

      port map(A => CO1_2, B => \framesync[2]_net_1\, Y => CO2_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \fsmdet_RNIIV9I[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmsync_ns_i_a3_0[6]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[1]_net_1\, 
        C => N_68, D => un70_fsmsta, Y => N_1007);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[0]_net_1\, B => seradr0apb(1), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_145_2, 
        Y => N_2171);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_3\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[27]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmsta[23]_net_1\, B => un1_fsmmod, C => 
        N_193, Y => N_166);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[2]_net_1\, B => seradr0apb(3), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_6, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    \serdat_RNIBFTA1[6]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[6]_net_1\, B => \sercon[6]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => \un1_rtn_4\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_1);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => \SDAInt\, B => N_108, C => N_126, D => 
        un136_framesync, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns\ : CFG4
      generic map(INIT => x"B888")

      port map(A => bsd7_tmp_6_am, B => bsd7_tmp_6_ns_1, C => 
        un92_fsmsta, D => CoreAPB3_0_APBmslave0_PWDATA(7), Y => 
        bsd7_tmp_6);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        C => un25_fsmsta_1, D => un135_ens1_7, Y => un25_fsmsta);
    
    \fsmmod_ns_0_a4_0[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => 
        N_1059_1, Y => N_1051);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \sersta_32_6[2]\, B => \sersta_32_7[2]\, C
         => N_23, D => \un1_fsmsta_2_1\, Y => \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, B => 
        \fsmmod[4]_net_1\, C => N_1040, D => un70_fsmsta, Y => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    un7_fsmsta_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[22]_net_1\, 
        Y => N_2178);
    
    PCLK_count1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"0405")

      port map(A => \sercon[7]_net_1\, B => ANC2, C => 
        \sercon[0]_net_1\, D => \PCLK_count1[3]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_1\);
    
    \fsmmod_ns_0[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_1064, B => N_1049, C => un115_fsmdet, D => 
        N_1048, Y => \fsmmod_ns[0]\);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_1\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_2181, B => \adrcompen\, C => N_26, Y => 
        fsmsta_8_28_307_a3_0_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => un1_fsmmod, B => SDAO_int_7_0_275_a5_0, C => 
        N_1466, D => SDAO_int_7_0_275_1, Y => N_1449);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \sercon[7]_net_1\, D => 
        \un1_pclk_count1_ov_1_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"003A")

      port map(A => \ack\, B => N_172, C => N_2177, D => 
        fsmsta_8_4_577_i_0, Y => N_2172_i_0);
    
    \fsmmod_ns_0_a4_0[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[1]_net_1\, B => \SCLSCL\, C => 
        \pedetect\, Y => N_1049);
    
    g0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => CONFIG_rega20_2);
    
    \fsmsta_RNO[25]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => N_172, B => N_2177, C => \fsmsta_8_i_0[25]\, 
        D => un136_framesync, Y => N_2175_i_0);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_6\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), Y => 
        un26_adrcompen_6);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync[2]_net_1\, D => \framesync[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[21]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1652, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_3_601_0_1);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns_1\ : CFG4
      generic map(INIT => x"1555")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_0_INT[0]\, 
        C => un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_ns_1);
    
    PCLK_count1_ov_1_sqmuxa_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[0]_net_1\, B => \sercon[1]_net_1\, Y
         => \PCLK_count1_ov_1_sqmuxa_0\);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => 
        un1_fsmmod, D => N_133, Y => N_2173_i_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_0_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \fsmmod_ns_i_a4_1_1[2]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \un151_framesync\, B => N_1035, C => 
        \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_i_a4_1_1[2]_net_1\);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \fsmmod_RNIJBT51[5]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmdet[3]_net_1\, Y => N_189);
    
    \un1_PCLK_count1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1_1_sqmuxa_1\, C => \PCLK_count1[1]_net_1\, Y
         => CO1);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[2]_net_1\, Y => N_76);
    
    \serdat_RNI59TA1[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_0_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \sercon_8[3]\, B => 
        CoreAPB3_0_APBmslave0_PWDATA(3), C => un5_penable_2, D
         => N_138, Y => \sercon_9[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[18]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.CO2\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, Y
         => CO2);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => \un1_rtn_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[21]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \fsmsta[21]_net_1\, B => N_2177, C => N_193, 
        Y => \fsmsta_s12[21]\);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    un7_fsmsta_i_0_o2_RNIFH161 : CFG3
      generic map(INIT => x"01")

      port map(A => N_2178, B => un57_fsmsta_1_0, C => 
        \un1_fsmsta_6\, Y => N_193);
    
    \sersta_RNIMKFQ1[4]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        seradr0apb(7), Y => N_1221);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \sercon[6]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_0_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"D555")

      port map(A => N_2176, B => N_2187, C => N_95, D => 
        \adrcomp_2_sqmuxa_i_a3_4\, Y => \adrcomp_2_sqmuxa_i_0\);
    
    \un2_framesync_1_1.CO1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CO0, B => \framesync[1]_net_1\, Y => CO1_2);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmmod[2]_net_1\, Y => SDAO_int_7_0_275_a5_0);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SDAO_int_RNITQ98 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_0_SDAO[0]\, Y => 
        COREI2C_0_0_SDAO_i(0));
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \COREI2C_0_0_SDAO[0]\, B => N_2177, C => 
        fsmsta_8_23_351_i_0_1, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \fsmsync_ns_0_a3_2_2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[4]_net_1\, Y
         => N_1002_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_9_509_0_1);
    
    \serCON_WRITE_PROC.sercon_8_0[3]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_161_2, B => N_163_2, C => \sercon_8_0_1[3]\, 
        D => \sercon_8_0_0[3]\, Y => \sercon_8[3]\);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"00BF")

      port map(A => \bsd7\, B => un57_fsmsta, C => 
        \un1_bsd7_1_sqmuxa[0]_net_1\, D => bsd7_9_iv_2, Y => 
        bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \indelay[1]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \fsmmod_ns_i_1[2]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => un70_fsmsta, B => 
        \fsmmod_ns_i_a4_1_1[2]_net_1\, C => \fsmmod[4]_net_1\, D
         => \fsmmod_ns_i_0[2]_net_1\, Y => 
        \fsmmod_ns_i_1[2]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_6[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[15]_net_1\, 
        C => \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_6[2]\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.ANC2\ : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, Y
         => ANC2);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(4), B => seradr0apb(2), C => 
        \serdat[3]_net_1\, D => \serdat[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_11_454_i_a6_2_0_0_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, Y => 
        N_2182);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_2, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"515F")

      port map(A => \fsmsta[11]_net_1\, B => N_2186, C => N_2177, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[1]_net_1\, C
         => \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2177, B => N_2178, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_0_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \fsmmod_ns_0_a4_0_1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \starto_en\, B => N_64, C => N_1040, D => 
        un115_fsmdet, Y => N_1059_1);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    un1_fsmsta_1_i_0_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[12]_net_1\, 
        C => \fsmsta[16]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => fsmsta_8_28_307, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => un135_ens1_7, B => \fsmsta[14]_net_1\, Y => 
        N_2196);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNIFFO81 : CFG4
      generic map(INIT => x"AF8C")

      port map(A => N_161_2, B => \pedetect\, C => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\, D => N_2181, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[0]\ : CFG4
      generic map(INIT => x"66F0")

      port map(A => \framesync[0]_net_1\, B => un8_nedetect, C
         => \framesync_7_m2[3]\, D => framesync_7_e2, Y => 
        \framesync_7[0]\);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_1[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1586_1, B => \sercon[6]_net_1\, Y => 
        N_163_2);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    PCLKint_ff_RNI9NL41 : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_0[3]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => \sercon[6]_net_1\, B => \COREI2C_0_0_INT[0]\, 
        C => N_1064, D => N_189, Y => \sercon_8_0_0[3]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \fsmsync_ns_i_0[6]\ : CFG4
      generic map(INIT => x"5C5F")

      port map(A => \SDAInt\, B => \COREI2C_0_0_INT[0]\, C => 
        \fsmsync[1]_net_1\, D => \sercon[4]_net_1\, Y => 
        \fsmsync_ns_i_0[6]_net_1\);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \un1_fsmsta_6\, B => un136_framesync, C => 
        \fsmsta_nxt_9_m_0[26]\, D => fsmsta_nxt_1_sqmuxa_18_s5_1, 
        Y => \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => \un1_fsmsta_6\, B => \fsmsta_nxt_9_m_0[21]\, 
        C => un136_framesync, D => \fsmsta_s12[21]\, Y => 
        \fsmsta_8[21]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_3_601_0_1, D => N_1717, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_ns_0_a4[5]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => \pedetect\, B => \SCLSCL\, C => un115_fsmdet, 
        D => \fsmmod[1]_net_1\, Y => N_1058);
    
    \serCON_WRITE_PROC.un5_penable_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => un5_penable_0);
    
    \fsmmod_ns_0_a4[0]\ : CFG4
      generic map(INIT => x"AAA2")

      port map(A => \fsmmod[6]_net_1\, B => \starto_en\, C => 
        N_1040, D => N_64, Y => N_1048);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sersta_RNIIGFQ1[3]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        seradr0apb(6), Y => N_1220);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"C5")

      port map(A => N_2196, B => \COREI2C_0_0_SDAO[0]\, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \ack\, B => N_2177, C => N_133, D => 
        fsmsta_8_28_307_a3_0_1, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \sersta_32_i_a2_7[3]\, D => \COREI2C_0_0_INT[0]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"1000")

      port map(A => \PCLK_count1_0_sqmuxa_2\, B => 
        \PCLK_count1_0_sqmuxa_1\, C => \PCLK_count1_1_sqmuxa_3\, 
        D => \PCLK_count1_1_sqmuxa_1\, Y => 
        \PCLK_count1_1_sqmuxa\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    serdat_2_sqmuxa : CFG4
      generic map(INIT => x"0020")

      port map(A => un92_fsmsta, B => un105_ens1, C => \pedetect\, 
        D => \COREI2C_0_0_INT[0]\, Y => \serdat_2_sqmuxa\);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[6]_net_1\, C
         => \fsmmod[1]_net_1\, Y => un16_fsmmod);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_RNITGHM\ : CFG3
      generic map(INIT => x"40")

      port map(A => \COREI2C_0_0_INT[0]\, B => un57_fsmsta, C => 
        \nedetect\, Y => bsd7_tmp_6_sn_m6_1);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"02")

      port map(A => N_2196, B => \COREI2C_0_0_SDAO[0]\, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        PCLK_count2_ov_6_1, C => CO1, D => \PCLK_count1_1_sqmuxa\, 
        Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[16]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_1[3]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        N_2177, D => N_2179, Y => N_162);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[12]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmmod_ns_i_o3_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_0_INT[0]\, B => \sercon[5]_net_1\, 
        Y => N_1035);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"00D0")

      port map(A => N_2186, B => N_2177, C => N_82, D => 
        un136_framesync, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \sersta_32_5[1]\, B => N_72_mux, C => 
        \sersta_32_4[1]\, Y => \sersta_32[1]\);
    
    \sersta_RNI64FQ1[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \fsmsync_ns_i_o3_0_i_o2[5]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_64, B => \fsmsync[5]_net_1\, Y => N_68);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[27]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_24_s4_1_0, Y => 
        \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG3
      generic map(INIT => x"54")

      port map(A => N_2181, B => fsmsta_8_5_555_a3_2, C => 
        fsmsta_8_5_555_a3_0_2, Y => fsmsta_8_5_555);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_0_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_0_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"7075")

      port map(A => \ack\, B => un13_adrcompen, C => 
        \adrcomp_2_sqmuxa_i_a2_1_5\, D => N_133, Y => N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    \serdat_RNIUIJ31[5]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(5), B => \serdat[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_0_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7[0]\ : CFG4
      generic map(INIT => x"07FF")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_e2_1, Y => 
        \framesync_7_m2[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => fsmsta_8_28_307);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    PCLK_count1_0_sqmuxa_4_1 : CFG3
      generic map(INIT => x"01")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \PCLK_count1_0_sqmuxa_4_1\);
    
    PCLK_count1_1_sqmuxa_1_0 : CFG4
      generic map(INIT => x"CCFA")

      port map(A => \sercon[1]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \sercon[7]_net_1\, D => 
        \PCLK_count1_1_sqmuxa_1_0_1\, Y => 
        \PCLK_count1_1_sqmuxa_1_0\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \fsmsta_RNO[19]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => un133_framesync, B => N_2199, C => N_157, D
         => N_2181, Y => N_2174_i_0);
    
    \serCON_WRITE_PROC.un5_penable_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => \un105_ens1_3\);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_0\ : CFG4
      generic map(INIT => x"CFEE")

      port map(A => N_2182, B => N_2181, C => \fsmsta[9]_net_1\, 
        D => N_2177, Y => fsmsta_8_4_577_i_0);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \COREI2C_0_0_INT[0]\, B => \fsmsta[9]_net_1\, 
        Y => \sersta_32_2[0]\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_0_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[4]_net_1\, Y => fsmsta_8_9_509_a4_0);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => fsmsta_8_20_379_i_0_a3_3, B => m7_3, C => 
        \fsmsta[1]_net_1\, D => \fsmsta[11]_net_1\, Y => N_72_mux);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \fsmsta[14]_net_1\, D => \fsmsta[12]_net_1\, Y => 
        un25_fsmsta_1);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFDC")

      port map(A => N_2177, B => un16_fsmmod, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_0_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO0, B => framesync_7_e2, C => 
        \framesync[1]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[1]\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => un16_fsmmod, B => \sercon_8_2[4]\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), D => un5_penable, Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => N_76, D => \fsmsync[4]_net_1\, Y => N_55_i_0);
    
    \FSMSTA_SYNC_PROC.un133_framesync\ : CFG3
      generic map(INIT => x"08")

      port map(A => un1_fsmmod, B => un91_ens1, C => 
        \fsmsta[23]_net_1\, Y => un133_framesync);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un133_framesync, B => N_2181, Y => 
        un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_1_sqmuxa_1\, D => 
        \PCLK_count1_1_sqmuxa\, Y => \PCLK_count1_10[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG4
      generic map(INIT => x"5554")

      port map(A => \fsmdet[3]_net_1\, B => un57_fsmsta_0, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un8_nedetect\ : CFG2
      generic map(INIT => x"E")

      port map(A => un70_fsmsta, B => \nedetect\, Y => 
        un8_nedetect);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    \un2_framesync_1_1.CO0\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \framesync[0]_net_1\, B => un70_fsmsta, C => 
        \nedetect\, Y => CO0);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    un1_fsmsta_2_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[24]_net_1\, B => \fsmsta[25]_net_1\, 
        Y => \un1_fsmsta_2_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"F7F5")

      port map(A => N_2178, B => \fsmsta[20]_net_1\, C => N_2188, 
        D => N_2177, Y => fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => \fsmmod[2]_net_1\, B => N_1064, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_138, B => un5_penable_2, Y => un5_penable);
    
    \serdat_RNIDHTA1[7]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[7]_net_1\, B => \sercon[7]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    PCLK_count1_0_sqmuxa_2 : CFG4
      generic map(INIT => x"0545")

      port map(A => \sercon[7]_net_1\, B => CO1_0, C => 
        \PCLK_count1[3]_net_1\, D => \PCLK_count1[2]_net_1\, Y
         => \PCLK_count1_0_sqmuxa_2\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1035, B => \sercon[4]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    PCLK_count1_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0070")

      port map(A => CO2, B => \PCLK_count1_0_sqmuxa_4_1\, C => 
        \PCLK_count1_1_sqmuxa_1_0\, D => \PCLK_count1_0_sqmuxa_3\, 
        Y => \PCLK_count1_1_sqmuxa_3\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => PCLK_count2_ov_6_0_a2_1_3, B => un16_fsmmod, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    un1_counter_rst_3 : CFG2
      generic map(INIT => x"B")

      port map(A => \PCLK_count1_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, Y => \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_0_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"ACAA")

      port map(A => \fsmsta[13]_net_1\, B => 
        \COREI2C_0_0_SDAO[0]\, C => N_2177, D => N_2196, Y => 
        N_82);
    
    \fsmsta_RNO[12]\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_124, B => N_2188, C => N_2186, Y => 
        N_1774_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_0_SDAO[0]\, Y => 
        N_172);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_3_0, B => 
        fsmsta_8_20_379_i_0_a3_3, C => N_2177, D => 
        fsmsta_8_20_379_i_0_a3_4, Y => N_145);
    
    adrcomp : SLE
      port map(D => N_2176, CLK => FAB_CCC_GL0, EN => 
        \adrcomp_2_sqmuxa_i_0\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG4
      generic map(INIT => x"1F10")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmdet[3]_net_1\, D => \fsmdet[1]_net_1\, Y => 
        N_1717);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[23]_net_1\, B => \fsmsta[7]_net_1\, Y
         => fsmsta_8_20_379_i_0_a3_3);
    
    un1_fsmsta_i_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[18]_net_1\, 
        Y => un135_ens1_7);
    
    \serCON_WRITE_PROC.un91_ens1_0_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \pedetect\, Y => un91_ens1);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \fsmsta[9]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => \fsmsta_cnst[0]\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \COREI2C_0_0_INT[0]\, B => un70_fsmsta, C => 
        \fsmmod[4]_net_1\, D => \sercon[4]_net_1\, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[26]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[8]_net_1\, B => \fsmsta[9]_net_1\, Y
         => N_145_2);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => fsmsta_8_5_555, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_68, B => \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \fsmmod[5]_net_1\, B => \nedetect\, C => 
        un115_fsmdet, D => N_1051, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_0_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \serCON_WRITE_PROC.un3_penable_1\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => \un3_penable_1\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => un57_fsmsta_0, D => un57_fsmsta_1_0, Y => 
        un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG2
      generic map(INIT => x"1")

      port map(A => fsmsta_8_2_647_i_0_0, B => N_2188, Y => 
        N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"70F0")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_pclk_count191\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_3\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[8]_net_1\, C
         => \fsmsta[2]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[22]\, B => un136_framesync, C
         => \fsmsta[22]_net_1\, D => N_2177, Y => \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => \un1_rtn_3\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_counter_rst_3\, D => 
        \PCLK_count1_1_sqmuxa_1\, Y => \PCLK_count1_10[1]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_4\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, Y => un135_ens1_4);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_64, D => N_1002_3, Y => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \bsd7_tmp\, B => \SCLInt\, C => 
        \COREI2C_0_0_INT[0]\, D => un57_fsmsta, Y => 
        bsd7_tmp_i_m_2);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"FFEA")

      port map(A => un105_ens1, B => \serdat_2_sqmuxa\, C => 
        \sercon[6]_net_1\, D => \serdat_1_sqmuxa_1\, Y => 
        \un1_serdat_2_sqmuxa\);
    
    \serdat_RNI7BTA1[4]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[4]_net_1\, B => \sercon[4]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[4]\);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \COREI2C_0_0_INT[0]\, B => N_1002, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_0_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_0_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"DCCC")

      port map(A => un105_ens1, B => \serdat_2_sqmuxa\, C => 
        \pedetect\, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_7\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[8]_net_1\, B => \fsmsta[7]_net_1\, C
         => un135_ens1_7, D => un135_ens1_4, Y => un135_ens1_7_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_26_328_a3_0_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => \fsmsta[23]_net_1\, B => \adrcomp\, Y => N_26);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[24]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \fsmsta[27]_net_1\, D => \fsmsta[26]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_3_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    SCLO_int_RNI7CA5 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_0_SCLO[0]\, Y => 
        COREI2C_0_0_SCLO_i(0));
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \fsmdet[1]_net_1\, B => fsmsta_8_3_601_a4_0, 
        C => N_1656, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_172, B => N_2182, C => N_2193, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, B => 
        N_1002_3, Y => N_1002);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_2\ : CFG4
      generic map(INIT => x"FF04")

      port map(A => \serdat[7]_net_1\, B => bsd7_tmp_6_sn_m6_1, C
         => un105_ens1, D => bsd7_9_iv_1, Y => bsd7_9_iv_2);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[27]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[3]_net_1\, B => \serdat[2]_net_1\, C
         => \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_0\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, C
         => \fsmsta[7]_net_1\, Y => un57_fsmsta_0);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[26]_net_1\, C => N_172, 
        Y => fsmsta_nxt_1_sqmuxa_18_s5_1);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ack\, B => \adrcompen\, C => N_2177, D => 
        N_26, Y => fsmsta_8_5_555_a3_0_2);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_0_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3340")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1586_1, Y => N_1624);
    
    adrcomp_2_sqmuxa_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[23]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => N_95);
    
    PCLK_count1_1_sqmuxa_1_0_1 : CFG4
      generic map(INIT => x"5008")

      port map(A => CO1_0, B => bclke, C => 
        \PCLK_count1[3]_net_1\, D => \PCLK_count1[2]_net_1\, Y
         => \PCLK_count1_1_sqmuxa_1_0_1\);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_0_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        \COREI2C_0_0_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_0_3\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[10]_net_1\, Y => fsmsta_8_3_601_a4_0);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    serdat_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \pedetect\, B => \sercon[6]_net_1\, C => 
        \un1_serdat40\, Y => \serdat_1_sqmuxa_1\);
    
    \fsmmod_RNO[4]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmmod_ns_i_1[2]_net_1\, B => un115_fsmdet, 
        C => N_1046, Y => N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \serDAT_WRITE_PROC.un105_ens1_0\ : CFG3
      generic map(INIT => x"10")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \un105_ens1_0\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_am\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \bsd7_tmp\, B => bsd7_tmp_6_sn_m6_1, C => 
        un105_ens1, Y => bsd7_tmp_6_am);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_1[3]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => un74_ens1, B => \adrcomp\, C => N_162, D => 
        N_163_2, Y => \sercon_8_0_1[3]\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2[7]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_2177, B => N_2181, C => \fsmsta[7]_net_1\, 
        D => N_172, Y => N_108);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_o3\ : CFG3
      generic map(INIT => x"FB")

      port map(A => N_1586_1, B => N_1656, C => \fsmsta_cnst[0]\, 
        Y => N_2188);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_0_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \fsmsta[29]_net_1\, B => \PCLKint_ff\, C => 
        \PCLKint\, D => \fsmsta[28]_net_1\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => N_1449, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_0_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[16]_net_1\, 
        C => \fsmsta[19]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_145, B => N_2181, C => N_166, D => 
        fsmsta_8_20_379_i_0_o2_0, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"3100")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_e2_1, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[6]_net_1\, B => \fsmsta[15]_net_1\, C
         => \fsmsta[2]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \CLK_COUNTER1_PROC.un12_pclk_count1_1.ANC1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, Y => CO1_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_9_509_0_1, D => N_1717, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_126, B => N_2181, C => un133_framesync, D
         => N_80, Y => N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"FBF8")

      port map(A => \PWDATA_i_m_1[7]\, B => un105_ens1, C => 
        \fsmdet[3]_net_1\, D => bsd7_tmp_i_m_2, Y => bsd7_9_iv_1);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG3
      generic map(INIT => x"04")

      port map(A => \fsmsta[29]_net_1\, B => N_145_2, C => 
        \fsmsta[25]_net_1\, Y => fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \fsmdet[1]_net_1\, B => fsmsta_8_9_509_a4_0, 
        C => N_1656, D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmmod_ns_0_a4_0_4[3]_net_1\, B => 
        un115_fsmdet, C => \fsmmod[3]_net_1\, D => N_1034, Y => 
        \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \sersta_32_2[0]\, B => N_72_mux, C => N_127, 
        D => \sersta_32_3[0]\, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        C => un135_ens1_7_0, D => un135_ens1_3, Y => un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0051")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp\, D => \fsmmod[0]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3[19]\ : CFG4
      generic map(INIT => x"0322")

      port map(A => un57_fsmsta_1_0, B => N_2177, C => \SDAInt\, 
        D => N_2178, Y => N_157);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \un3_penable_1\, B => N_138, C => 
        \un105_ens1_0\, D => \un105_ens1_3\, Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    \fsmsync_ns_i_a3_1_0_a2_2[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[3]_net_1\, C
         => \fsmmod[1]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_0_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \sersta_RNIA8FQ1[1]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[4]\, C => \sersta[1]_net_1\, D => 
        seradr0apb(4), Y => N_1218);
    
    \fsmsync_RNO[1]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_1007, B => \fsmsync_ns_i_0[6]_net_1\, C => 
        N_1002, Y => N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1058, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_0_INT[0]\, 
        C => \fsmsta[24]_net_1\, D => \fsmsta[28]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_0_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[3]\ : CFG4
      generic map(INIT => x"7D28")

      port map(A => framesync_7_e2, B => CO2_0, C => 
        \framesync[3]_net_1\, D => \framesync_7_m2[3]\, Y => 
        \framesync_7[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    PCLK_count1_1_sqmuxa_1 : CFG4
      generic map(INIT => x"8CCC")

      port map(A => bclke, B => PCLK_count2_ov_6_1, C => 
        \sercon[7]_net_1\, D => \PCLK_count1_ov_1_sqmuxa_0\, Y
         => \PCLK_count1_1_sqmuxa_1\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[5]_net_1\, B => \fsmsync[2]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG4
      generic map(INIT => x"0307")

      port map(A => \fsmmod[0]_net_1\, B => \nedetect\, C => 
        \fsmmod[4]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \fsmmod_ns_i_0[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_1586_1, B => \fsmsta[8]_net_1\, C => N_2177, 
        D => N_172, Y => fsmsta_8_5_555_a3_2);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => \un1_rtn_3\);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    
    \sersta_RNIECFQ1[2]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        \sercon[5]_net_1\, Y => N_1219);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmdet[3]_net_1\, B => un139_ens1_0, C => 
        \fsmdet[1]_net_1\, Y => framesync_7_e2_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C is

    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          COREI2C_0_0_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          un3_penable                                : in    std_logic;
          bclke                                      : out   std_logic;
          un561_psel_4                               : out   std_logic;
          CONFIG_rega20_2                            : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_0_SDA_IO_Y                 : in    std_logic;
          un105_ens1_3                               : out   std_logic;
          BIBUF_COREI2C_0_0_SCL_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          un3_penable_1                              : out   std_logic;
          un5_penable_0                              : out   std_logic;
          un105_ens1_0                               : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_138                                      : in    std_logic;
          un5_penable_2                              : in    std_logic
        );

end COREI2C;

architecture DEF_ARCH of COREI2C is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6
    port( COREI2C_0_0_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0) := (others => 'U');
          seradr0apb                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          CONFIG_rega20_2                            : out   std_logic;
          bclke                                      : in    std_logic := 'U';
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_0_SDA_IO_Y                 : in    std_logic := 'U';
          un105_ens1_3                               : out   std_logic;
          BIBUF_COREI2C_0_0_SCL_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          un3_penable_1                              : out   std_logic;
          un5_penable_0                              : out   std_logic;
          un105_ens1_0                               : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_138                                      : in    std_logic := 'U';
          un5_penable_2                              : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\, \bclk_ff\, \bclk_ff0\, bclke_net_1
         : std_logic;

    for all : COREI2CREAL_6
	Use entity work.COREI2CREAL_6(DEF_ARCH);
begin 

    bclke <= bclke_net_1;

    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \serADR0_WRITE_PROCa.un3_penable_4\ : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(1), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => un561_psel_4);
    
    \bclke\ : CFG2
      generic map(INIT => x"2")

      port map(A => \bclk_ff0\, B => \bclk_ff\, Y => bclke_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    bclk_ff0 : SLE
      port map(D => FAB_CCC_GL0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bclk_ff0\);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    bclk_ff : SLE
      port map(D => \bclk_ff0\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bclk_ff\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6
      port map(COREI2C_0_0_SDAO_i(0) => COREI2C_0_0_SDAO_i(0), 
        COREI2C_0_0_SCLO_i(0) => COREI2C_0_0_SCLO_i(0), 
        COREI2C_0_0_INT(0) => COREI2C_0_0_INT(0), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, CONFIG_rega20_2 => 
        CONFIG_rega20_2, bclke => bclke_net_1, N_1221 => N_1221, 
        N_1217 => N_1217, N_1220 => N_1220, N_1218 => N_1218, 
        N_1219 => N_1219, BIBUF_COREI2C_0_0_SDA_IO_Y => 
        BIBUF_COREI2C_0_0_SDA_IO_Y, un105_ens1_3 => un105_ens1_3, 
        BIBUF_COREI2C_0_0_SCL_IO_Y => BIBUF_COREI2C_0_0_SCL_IO_Y, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, un3_penable_1 => 
        un3_penable_1, un5_penable_0 => un5_penable_0, 
        un105_ens1_0 => un105_ens1_0, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, N_138 => N_138, 
        un5_penable_2 => un5_penable_2);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( MSS_READY                                : out   std_logic;
          FAB_CCC_GL0                              : in    std_logic;
          POWER_ON_RESET_N                         : in    std_logic;
          M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \POWER_ON_RESET_N_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \POWER_ON_RESET_N_q1\, \RESET_N_M2F_q1\, 
        \FIC_2_APB_M_PRESET_N_q1\, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \MSS_HPMS_READY_int_3\
         : std_logic;

begin 


    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => POWER_ON_RESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \POWER_ON_RESET_N_clk_base\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_q1\);
    
    MSS_HPMS_READY_int_RNILPQ3 : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => \POWER_ON_RESET_N_clk_base\, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_0 is

    port( COREI2C_0_1_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0);
          seradr0apb                                 : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_1_SCL_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_1_SDA_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          un3_penable_1                              : out   std_logic;
          un105_ens1_3                               : in    std_logic;
          un105_ens1_1                               : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic;
          un5_penable_1                              : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          bclke                                      : in    std_logic;
          N_138                                      : in    std_logic
        );

end COREI2CREAL_6_0;

architecture DEF_ARCH of COREI2CREAL_6_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_1_SDAO[0]\, \COREI2C_0_1_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_1_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        un1_serdat_2_sqmuxa_0, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, N_1665, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, N_1470, \ack\, ack_7, N_1449, 
        SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, bsd7_tmp_6, \bsd7\, 
        bsd7_9_iv_i_0, \adrcomp\, \adrcomp_2_sqmuxa_i_0_0_i\, 
        adrcomp_2_sqmuxa_i_0_0, \PCLKint\, PCLKint_3, 
        un1_pclkint4_i_0, \ack_bit\, \ack_bit_1_sqmuxa\, 
        \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_0, un1_rtn_3_0, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, PCLK_count2_ov_6_1, 
        \PCLK_count1_1_sqmuxa_1\, CO1, N_1586_1, un133_framesync, 
        \fsmsta_cnst[0]\, un136_framesync, N_997, un70_fsmsta, 
        N_1046, \adrcomp_2_sqmuxa_i_a3_2_0\, N_1622_2, 
        \adrcomp_2_sqmuxa_i_o2_1_3\, \sersta_32_5[2]\, N_66, N_84, 
        N_2177, N_2181, N_2173_i_1, N_133, un1_fsmmod, N_36_i_1, 
        N_2196, N_2186, \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, 
        fsmsta_8_3_601_0_1, N_1717, fsmsta_8_3_601_0, N_1652, 
        fsmsta_8_9_509_0_1, fsmsta_8_9_509_0, 
        \adrcomp_2_sqmuxa_i_a2_1_2\, un13_adrcompen, 
        \adrcomp_2_sqmuxa_i_a2_1_1_0\, N_168, 
        \adrcomp_2_sqmuxa_i_a2_1_1\, \adrcomp_2_sqmuxa_i_a2_1_0\, 
        CO2, \PCLK_count1_1_sqmuxa_2_1\, \PCLK_count1_1_sqmuxa_2\, 
        \un1_pclk_count1_ov_1_1\, \un1_pclk_count1_ov_1\, 
        \PCLK_count1_1_sqmuxa_0_1_0\, \PCLK_count1_1_sqmuxa_0\, 
        \PRDATA_3_1_1[7]\, \PRDATA_3_1_1[3]\, \PRDATA_3_1[4]\, 
        \PRDATA_3_1_1[6]\, \PRDATA_3_1_1[5]\, \fsmsta_8_ns_1[28]\, 
        \fsmsta_8_ns_1[29]\, \fsmsta_8_ns_1[18]\, 
        \fsmsta_8_ns_1[16]\, bsd7_tmp_6_ns_1, bsd7_tmp_6_am_1, 
        un105_ens1, un57_fsmsta, N_2179, N_161_2, N_2171, 
        \fsmsta_8_0_a2_1[7]\, fsmsta_8_5_555_a3_0_2, 
        fsmsta_8_5_555_a3_2, N_2193, \un1_fsmsta_6\, N_2199, 
        bsd7_tmp_6_sn_m6_0, PCLK_count2_ov_6_0_a2_1_0, 
        \sersta_32_2[0]\, un111_fsmdet_0, \sersta_32_i_a2_5[3]\, 
        \PCLK_count1_ov_1_sqmuxa_0\, \adrcomp_2_sqmuxa_i_a3_2\, 
        N_629, un139_ens1_0, fsmsta_8_20_379_i_0_a3_3, 
        \adrcomp_2_sqmuxa_i_o2_1_1\, \un1_fsmsta_1_i_0_o2_0\, 
        N_127, N_23, N_64, un135_ens1_2, N_67, un10_sclscl, 
        N_1002_3, N_2178, N_26, N_145_2, \un151_framesync\, 
        N_1196, N_1197, N_1198, \serdat_i_m_1[7]\, bsd7_tmp_i_m_1, 
        SDAO_int_7_0_275_1, SDAO_int_7_0_275_a5_0, un141_ens1_2, 
        fsmsta_8_28_307_a3_0_0, \SDAO_int_1_sqmuxa_3\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_10_476_i_a6_1, 
        \sersta_32_5[1]\, \sersta_32_4[1]\, \sersta_32_3[0]\, 
        \fsmmod_ns_i_a4_1_0[2]_net_1\, fsmsta_8_20_379_i_0_a3_4, 
        fsmsta_8_20_379_i_0_a3_3_0, \sersta_32_i_a2_7[4]\, 
        \sersta_32_i_a2_6[4]\, \sersta_32_4[2]\, un135_ens1_5, 
        un135_ens1_4, un135_ens1_3, fsmsta_nxt_1_sqmuxa_24_s4_1_0, 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0, un25_fsmsta_1, 
        \sersta_32_i_a2_8[3]\, \sersta_32_i_a2_7[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, m7_3, 
        un13_adrcompen_4, N_1064, un33_fsmsta, \un3_penable_1\, 
        framesync_7_sm0, PCLK_count2_ov_6_0_a2_1_4_tz, N_1034, 
        un16_fsmmod, N_1040, N_76, \un1_pclk_count1_ov\, CO1_0, 
        CO1_1, \adrcomp_2_sqmuxa_i_a3_3\, 
        \fsmmod_ns_i_0[2]_net_1\, fsmsta_8_10_476_i_0, 
        \SDAO_int_1_sqmuxa_4\, PCLK_count2_ov_6_0_a2_1_3, 
        \adrcomp_2_sqmuxa_i_0_0_0\, \sercon_8_2[4]\, 
        \sersta_32_i_a2_9[4]\, \sersta_32_7[2]\, 
        \sersta_32_i_a2_10[3]\, N_2192, N_72_mux, N_104, N_1044, 
        un19_framesync, un25_fsmsta, un25_framesync, N_1002, 
        \un105_ens1_1\, \un5_penable_1\, N_130, N_995, un74_ens1, 
        N_63, \un1_pclk_count191\, N_1732, CO2_0, N_1656, N_1041, 
        N_154, N_191, N_155, N_120, N_121, N_124, 
        \adrcomp_2_sqmuxa_i_a3_4\, \SDAO_int_1_sqmuxa_7\, 
        \fsmsync_ns_i_1[6]_net_1\, framesync_7_e2, N_1054, 
        un115_fsmdet, \fsmsta_nxt_9_m[22]\, un135_ens1, N_163, 
        N_162, \fsmsta_nxt_9_m[27]\, \fsmsta_nxt_9_m[26]\, 
        \fsmsta_nxt_9_m[21]\, N_157, N_165, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, N_1060, N_70, 
        \PCLK_count1_0_sqmuxa_3\, N_1624, N_160, N_1727_2, N_126, 
        \fsmsta_8_i_0[25]\, N_80, N_82, 
        \PCLK_count1_1_sqmuxa_1_0\, \fsmmod_ns_0_0[0]_net_1\, 
        fsmsta_8_20_379_i_0_o2_0, \fsmsync_ns_0_0_1[0]_net_1\, 
        fsmsta_8_23_351_i_0_1, \un1_ens1_pre_1_sqmuxa_0_a2_1\, 
        N_1465, N_166, N_145, \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        N_86, un92_fsmsta, un1_fsmsta_10_i_0, 
        \serdat_2_sqmuxa_1_0\, \PWDATA_i_m_1[7]\, 
        \sercon_8_0_2[3]\, fsmsta_8_2_647_i_0_0, N_1059, N_1051, 
        N_1486, \serdat_0_sqmuxa\, un134_fsmsta, 
        \framesync_7_m2[3]\, N_161, N_1466, N_152, bsd7_9_iv_1, 
        \un1_serdat40\, \un1_bsd7_1_sqmuxa[0]_net_1\, bsd7_9_iv_2, 
        \serdat_1_sqmuxa_1\, \un1_counter_rst_3\, 
        \un1_serdat_2_sqmuxa_1\ : std_logic;

begin 

    COREI2C_0_1_INT(0) <= \COREI2C_0_1_INT[0]\;
    un3_penable_1 <= \un3_penable_1\;
    un105_ens1_1 <= \un105_ens1_1\;
    un5_penable_1 <= \un5_penable_1\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \un151_framesync\, B => N_2177, C => N_191, Y
         => un1_fsmsta_10_i_0);
    
    \un1_bsd7_1_sqmuxa[0]\ : CFG3
      generic map(INIT => x"A1")

      port map(A => un105_ens1, B => \nedetect\, C => 
        \COREI2C_0_1_INT[0]\, Y => \un1_bsd7_1_sqmuxa[0]_net_1\);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    \un2_framesync_1_1.CO2\ : CFG2
      generic map(INIT => x"8")

      port map(A => CO1_1, B => \framesync[2]_net_1\, Y => CO2_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_0_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_26, B => \adrcompen\, Y => 
        fsmsta_8_28_307_a3_0_0);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_145_2, 
        Y => N_2171);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_3\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[19]_net_1\, 
        C => \fsmsta[4]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_191, B => \un1_fsmsta_6\, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => N_166);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_0);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    SDAO_int_RNIUE82 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_1_SDAO[0]\, Y => 
        COREI2C_0_1_SDAO_i(0));
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns\ : CFG4
      generic map(INIT => x"5404")

      port map(A => \fsmdet[3]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => bsd7_tmp_6_ns_1, D
         => bsd7_tmp_6_am_1, Y => bsd7_tmp_6);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => un25_fsmsta_1, 
        C => \fsmsta[18]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        un25_fsmsta);
    
    \fsmmod_ns_0_a4_0[1]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => N_1044, 
        D => un115_fsmdet, Y => N_1051);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sersta_32_5[2]\, B => \sersta_32_7[2]\, C
         => un135_ens1_2, D => \un1_fsmsta_1_i_0_o2_0\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1041, B => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, 
        C => N_1040, Y => \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    un7_fsmsta_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[22]_net_1\, 
        Y => N_2178);
    
    \fsmmod_ns_0[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un115_fsmdet, B => \fsmmod_ns_0_0[0]_net_1\, 
        C => N_1064, Y => \fsmmod_ns[0]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    \fsmmod_ns_0_0[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => N_1044, D => un10_sclscl, Y => 
        \fsmmod_ns_0_0[0]_net_1\);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    adrcomp_2_sqmuxa_i_a2_1_1 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(7), B => seradr0apb(4), C => 
        \serdat[6]_net_1\, D => \serdat[3]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_1\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => un1_fsmmod, B => SDAO_int_7_0_275_1, C => 
        SDAO_int_7_0_275_a5_0, D => N_1466, Y => N_1449);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_am_RNO\ : CFG2
      generic map(INIT => x"4")

      port map(A => \COREI2C_0_1_INT[0]\, B => \nedetect\, Y => 
        bsd7_tmp_6_sn_m6_0);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CEFF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \un1_pclk_count1_ov_1_1\, D => 
        \sercon[7]_net_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => un139_ens1_0, Y => 
        framesync_7_sm0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_2181, B => N_121, C => N_154, D => N_155, Y
         => N_2172_i_0);
    
    adrcomp_2_sqmuxa_i_0_0_i : CFG3
      generic map(INIT => x"15")

      port map(A => \adrcomp_2_sqmuxa_i_0_0_0\, B => 
        \COREI2C_0_1_INT[0]\, C => N_2192, Y => 
        \adrcomp_2_sqmuxa_i_0_0_i\);
    
    \fsmsta_RNO[25]\ : CFG3
      generic map(INIT => x"01")

      port map(A => un136_framesync, B => N_154, C => 
        \fsmsta_8_i_0[25]\, Y => N_2175_i_0);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_2_0\, Y
         => \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \fsmsta[17]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_2[3]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \sercon[6]_net_1\, B => \adrcomp\, C => 
        N_1586_1, D => un74_ens1, Y => N_163);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1652, D => un1_fsmmod, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_3_601_0_1);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_ns_1\ : CFG3
      generic map(INIT => x"7F")

      port map(A => un105_ens1, B => \COREI2C_0_1_INT[0]\, C => 
        un57_fsmsta, Y => bsd7_tmp_6_ns_1);
    
    PCLK_count1_ov_1_sqmuxa_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[0]_net_1\, B => \sercon[1]_net_1\, Y
         => \PCLK_count1_ov_1_sqmuxa_0\);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_1_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        N_161_2, Y => N_161);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \un1_PCLK_count1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1_1_sqmuxa_1\, C => \PCLK_count1[1]_net_1\, Y
         => CO1);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_66, B => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"FE0E")

      port map(A => \sercon_8_0_2[3]\, B => N_161, C => 
        un5_penable, D => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \sercon_9[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[18]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2171, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    adrcomp_2_sqmuxa_i_a2_1 : CFG4
      generic map(INIT => x"002A")

      port map(A => \adrcomp_2_sqmuxa_i_a2_1_2\, B => \ack\, C
         => un13_adrcompen, D => \adrcomp_2_sqmuxa_i_a2_1_1_0\, Y
         => N_168);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \sercon[6]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_1_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \COREI2C_0_1_INT[0]\, B => N_2192, C => 
        \adrcomp_2_sqmuxa_i_0_0_0\, D => N_152, Y => 
        adrcomp_2_sqmuxa_i_0_0);
    
    \un2_framesync_1_1.CO1\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp_2_sqmuxa_i_a3_2\, B => 
        \framesync[1]_net_1\, Y => CO1_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_629, B => \fsmmod[2]_net_1\, Y => 
        SDAO_int_7_0_275_a5_0);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_2181, B => fsmsta_8_23_351_i_0_1, C => 
        N_1656, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \fsmsync_ns_0_a3_2_2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[4]_net_1\, Y
         => N_1002_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_9_509_0_1);
    
    \sersta_RNIMT2J1[3]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        seradr0apb(6), Y => N_1220);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0D0F")

      port map(A => un92_fsmsta, B => \bsd7\, C => bsd7_9_iv_2, D
         => \un1_bsd7_1_sqmuxa[0]_net_1\, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[0]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_RNI20H61[5]\ : CFG4
      generic map(INIT => x"FEF0")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmsta_cnst[0]\, D => \fsmdet[3]_net_1\, Y => 
        N_1622_2);
    
    \serdat_RNIDP2S[6]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[6]_net_1\, B => \sercon[6]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \serSTA_WRITE_PROC.sersta_32_5[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[24]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_5[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_2177, B => N_172, Y => N_154);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(3), B => seradr0apb(2), C => 
        \serdat[2]_net_1\, D => \serdat[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a3_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta_cnst[0]\, B => \fsmdet[3]_net_1\, Y
         => N_1732);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    adrcomp_2_sqmuxa_i_a3 : CFG4
      generic map(INIT => x"F010")

      port map(A => N_133, B => \ack\, C => 
        \adrcomp_2_sqmuxa_i_a3_4\, D => N_168, Y => N_152);
    
    \serCON_WRITE_PROC.sercon_8_0_a3[3]\ : CFG4
      generic map(INIT => x"CC08")

      port map(A => \fsmdet[3]_net_1\, B => \sercon[6]_net_1\, C
         => N_629, D => N_1064, Y => N_160);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_1, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"4577")

      port map(A => \fsmsta[11]_net_1\, B => N_2177, C => N_2186, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[1]_net_1\, C
         => \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    adrcomp_2_sqmuxa_i_0_0_0 : CFG2
      generic map(INIT => x"E")

      port map(A => un16_fsmmod, B => N_1586_1, Y => 
        \adrcomp_2_sqmuxa_i_0_0_0\);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2177, B => N_2178, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, Y
         => N_629);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_1_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    adrcomp_2_sqmuxa_i_a3_2 : CFG2
      generic map(INIT => x"8")

      port map(A => \framesync[0]_net_1\, B => \nedetect\, Y => 
        \adrcomp_2_sqmuxa_i_a3_2\);
    
    un1_fsmsta_1_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => 
        \fsmsta[12]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => N_1470, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[14]_net_1\, 
        C => \fsmsta[18]_net_1\, Y => N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[0]\ : CFG4
      generic map(INIT => x"66F0")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync_7_m2[3]\, D => framesync_7_e2, Y => 
        \framesync_7[0]\);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[26]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_18_s5_1_0, Y => 
        \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \CLK_COUNTER1_PROC.un1_bclke_1.CO2\ : CFG3
      generic map(INIT => x"01")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[21]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \serdat_RNIUJ1R[4]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(4), B => \serdat[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_3_601_0_1, D => N_1717, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    PCLK_count1_1_sqmuxa_0 : CFG4
      generic map(INIT => x"FAFE")

      port map(A => \sercon[1]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \sercon[7]_net_1\, D => 
        \PCLK_count1_1_sqmuxa_0_1_0\, Y => 
        \PCLK_count1_1_sqmuxa_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \sersta_RNIAH2J1[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_m2\ : CFG4
      generic map(INIT => x"C5C0")

      port map(A => \fsmsta[23]_net_1\, B => \fsmsta[9]_net_1\, C
         => N_2177, D => un1_fsmmod, Y => N_121);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \COREI2C_0_1_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_155, B => fsmsta_8_28_307_a3_0_0, C => 
        N_133, D => N_2181, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \sersta_32_i_a2_7[3]\, D => \COREI2C_0_1_INT[0]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    un1_fsmsta_1_i_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        Y => \un1_fsmsta_1_i_0_o2_0\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \PCLK_count1_1_sqmuxa_1_0\, B => 
        \PCLK_count1_1_sqmuxa_1\, C => \PCLK_count1_1_sqmuxa_2\, 
        D => \PCLK_count1_1_sqmuxa_0\, Y => 
        \PCLK_count1_1_sqmuxa\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[6]_net_1\, C
         => \fsmmod[1]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_1_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_36_i_1);
    
    PCLKint_ff_RNICLRM : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        PCLK_count2_ov_6_1, C => CO1, D => \PCLK_count1_1_sqmuxa\, 
        Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[16]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_2177, B => \ack\, Y => N_155);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    adrcomp_2_sqmuxa_i_a2_1_1_0 : CFG4
      generic map(INIT => x"6FFF")

      port map(A => seradr0apb(1), B => \serdat[0]_net_1\, C => 
        \adrcomp_2_sqmuxa_i_a2_1_1\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_1_0\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_1[3]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        N_2177, D => N_2179, Y => N_162);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \serdat_RNI0M1R[5]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(5), B => \serdat[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => N_2186, B => N_2177, C => un136_framesync, D
         => N_82, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \sersta_32_5[1]\, B => N_72_mux, C => 
        \sersta_32_4[1]\, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[27]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_24_s4_1_0, Y => 
        \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG3
      generic map(INIT => x"54")

      port map(A => N_2181, B => fsmsta_8_5_555_a3_0_2, C => 
        fsmsta_8_5_555_a3_2, Y => N_1665);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_1_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_1_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_1_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7[0]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_m2[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => N_1470);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNIJJUR : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        un136_framesync, C => \pedetect\, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    PCLK_count1_1_sqmuxa_1_0 : CFG4
      generic map(INIT => x"00BF")

      port map(A => \PCLK_count1[3]_net_1\, B => CO2, C => bclke, 
        D => \PCLK_count1_0_sqmuxa_3\, Y => 
        \PCLK_count1_1_sqmuxa_1_0\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    PCLK_count1_1_sqmuxa_2 : CFG4
      generic map(INIT => x"CCCE")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \sercon[7]_net_1\, C => CO2, D => 
        \PCLK_count1_1_sqmuxa_2_1\, Y => \PCLK_count1_1_sqmuxa_2\);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \serdat_RNI7J2S[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_1_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \fsmsta_RNO[19]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_2199, B => un136_framesync, C => N_157, Y
         => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \COREI2C_0_1_INT[0]\, B => \sercon[5]_net_1\, 
        C => N_1041, D => \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => 
        N_1054);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \COREI2C_0_1_INT[0]\, B => \fsmsta[9]_net_1\, 
        Y => \sersta_32_2[0]\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => m7_3, B => fsmsta_8_20_379_i_0_a3_3, C => 
        \fsmsta[1]_net_1\, D => \fsmsta[11]_net_1\, Y => N_72_mux);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \fsmsta[14]_net_1\, D => \fsmsta[12]_net_1\, Y => 
        un25_fsmsta_1);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFDC")

      port map(A => N_2177, B => un16_fsmmod, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_1_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"3ACA")

      port map(A => \fsmdet[3]_net_1\, B => \framesync[1]_net_1\, 
        C => framesync_7_e2, D => \adrcomp_2_sqmuxa_i_a3_2\, Y
         => \framesync_7[1]\);
    
    serdat_2_sqmuxa_1_0 : CFG4
      generic map(INIT => x"0040")

      port map(A => \COREI2C_0_1_INT[0]\, B => un57_fsmsta, C => 
        \pedetect\, D => \fsmdet[3]_net_1\, Y => 
        \serdat_2_sqmuxa_1_0\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => un16_fsmmod, B => \sercon_8_2[4]\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), D => un5_penable, Y => 
        \sercon_9[4]\);
    
    \sersta_RNIEL2J1[1]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1[4]\, C => \sersta[1]_net_1\, D => 
        \sercon[4]_net_1\, Y => N_1218);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_76, Y => N_55_i_0);
    
    \FSMSTA_SYNC_PROC.un133_framesync\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \pedetect\, B => \fsmsta[23]_net_1\, C => 
        un1_fsmmod, D => N_2177, Y => un133_framesync);
    
    \sersta_RNIIP2J1[2]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        \sercon[5]_net_1\, Y => N_1219);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG3
      generic map(INIT => x"FE")

      port map(A => N_1586_1, B => un133_framesync, C => 
        \fsmsta_cnst[0]\, Y => un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_1_sqmuxa_1\, D => 
        \PCLK_count1_1_sqmuxa\, Y => \PCLK_count1_10[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, Y => 
        un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG3
      generic map(INIT => x"37")

      port map(A => N_67, B => \fsmsync[4]_net_1\, C => N_66, Y
         => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \serDAT_WRITE_PROC.un105_ens1_1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => un105_ens1_3, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \un105_ens1_1\);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"3AFF")

      port map(A => \COREI2C_0_1_SDAO[0]\, B => 
        \fsmsta[20]_net_1\, C => N_2177, D => N_2178, Y => 
        fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => \fsmmod[2]_net_1\, B => N_1064, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG3
      generic map(INIT => x"80")

      port map(A => \un3_penable_1\, B => \un5_penable_1\, C => 
        N_138, Y => un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_1_INT[0]\, 
        C => \sercon[5]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => PCLK_count2_ov_6_0_a2_1_3, B => un16_fsmmod, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    un1_counter_rst_3 : CFG2
      generic map(INIT => x"B")

      port map(A => \PCLK_count1_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, Y => \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_1_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"CACC")

      port map(A => \COREI2C_0_1_SDAO[0]\, B => 
        \fsmsta[13]_net_1\, C => N_2177, D => N_2196, Y => N_82);
    
    \fsmsta_RNO[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1656, B => N_2186, C => N_2181, D => N_124, 
        Y => N_1774_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_1_SDAO[0]\, Y => 
        N_172);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_3_0, B => 
        fsmsta_8_20_379_i_0_a3_3, C => N_2177, D => 
        fsmsta_8_20_379_i_0_a3_4, Y => N_145);
    
    adrcomp : SLE
      port map(D => \adrcomp_2_sqmuxa_i_0_0_i\, CLK => 
        FAB_CCC_GL0, EN => adrcomp_2_sqmuxa_i_0_0, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \adrcomp\);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \fsmdet[3]_net_1\, B => N_629, C => 
        \fsmdet[1]_net_1\, Y => N_1717);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_5\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => un135_ens1_2, Y => un135_ens1_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[23]_net_1\, B => \fsmsta[7]_net_1\, Y
         => fsmsta_8_20_379_i_0_a3_3);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \fsmsta[9]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => \fsmsta_cnst[0]\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0_RNIFLPL\ : CFG2
      generic map(INIT => x"1")

      port map(A => un57_fsmsta_1_0, B => N_2178, Y => N_191);
    
    \fsmmod_ns_i_o3[2]\ : CFG3
      generic map(INIT => x"BF")

      port map(A => N_997, B => un70_fsmsta, C => 
        \fsmmod[4]_net_1\, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[26]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, Y
         => N_145_2);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => N_1665, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \fsmsync[5]_net_1\, B => N_64, C => 
        \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \fsmmod[5]_net_1\, B => \nedetect\, C => 
        un115_fsmdet, D => N_1051, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_1_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \serCON_WRITE_PROC.un3_penable_1\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => \un3_penable_1\);
    
    PCLK_count1_1_sqmuxa_0_1_0 : CFG4
      generic map(INIT => x"377F")

      port map(A => \sercon[0]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => 
        \PCLK_count1_1_sqmuxa_0_1_0\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => un135_ens1_2, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_2181, B => fsmsta_8_2_647_i_0_0, C => 
        N_1656, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \fsmsta[23]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp_2_sqmuxa_i_a3_3\, D => \fsmmod[1]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[20]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[22]\, B => un136_framesync, C
         => \fsmsta[22]_net_1\, D => N_2177, Y => \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_counter_rst_3\, D => 
        \PCLK_count1_1_sqmuxa_1\, Y => \PCLK_count1_10[1]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_4\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, Y => un135_ens1_4);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_64, D => N_1002_3, Y => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SCLInt\, B => \COREI2C_0_1_INT[0]\, C => 
        \bsd7_tmp\, Y => bsd7_tmp_i_m_1);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \serdat_2_sqmuxa_1_0\, B => \sercon[6]_net_1\, 
        C => un105_ens1, D => \serdat_1_sqmuxa_1\, Y => 
        un1_serdat_2_sqmuxa_0);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \indelay[1]_net_1\, B => \indelay[3]_net_1\, 
        Y => N_66);
    
    \sersta_RNIQ13J1[4]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        seradr0apb(7), Y => N_1221);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1002, B => \COREI2C_0_1_INT[0]\, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_1_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FF7F")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_66, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_1_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"0E0A")

      port map(A => \serdat_2_sqmuxa_1_0\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_26_328_a3_0_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => \fsmsta[23]_net_1\, B => \adrcomp\, Y => N_26);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    SCLO_int_RNI809F : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_1_SCLO[0]\, Y => 
        COREI2C_0_1_SCLO_i(0));
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \serdat_RNIFR2S[7]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[7]_net_1\, B => \sercon[7]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_3_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    PCLK_count1_1_sqmuxa_2_1 : CFG4
      generic map(INIT => x"0111")

      port map(A => \sercon[0]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => 
        \PCLK_count1_1_sqmuxa_2_1\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[10]_net_1\, C => 
        N_1727_2, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, C => 
        N_2193, D => N_172, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, B => 
        N_1002_3, Y => N_1002);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_2\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => \fsmdet[3]_net_1\, B => \PWDATA_i_m_1[7]\, C
         => un105_ens1, D => bsd7_9_iv_1, Y => bsd7_9_iv_2);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_2_RNO\ : CFG4
      generic map(INIT => x"0002")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => \fsmdet[3]_net_1\, 
        D => \COREI2C_0_1_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[27]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[3]_net_1\, B => \serdat[2]_net_1\, C
         => \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[26]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ack\, B => \adrcompen\, C => N_2177, D => 
        N_26, Y => fsmsta_8_5_555_a3_0_2);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_1_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3430")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1586_1, D => un1_fsmmod, Y => N_1624);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_1_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => \nedetect\, B => \COREI2C_0_1_INT[0]\, C => 
        \serdat[7]_net_1\, Y => \serdat_i_m_1[7]\);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    serdat_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \pedetect\, B => \sercon[6]_net_1\, C => 
        \un1_serdat40\, Y => \serdat_1_sqmuxa_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_1046, B => \fsmmod_ns_i_0[2]_net_1\, C => 
        N_1054, D => un115_fsmdet, Y => N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_am\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => un57_fsmsta, B => un105_ens1, C => \bsd7_tmp\, 
        D => bsd7_tmp_6_sn_m6_0, Y => bsd7_tmp_6_am_1);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \serCON_WRITE_PROC.un5_penable_1\ : CFG4
      generic map(INIT => x"0004")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(0), B => 
        CONFIG_rega20_2, C => CoreAPB3_0_APBmslave0_PADDR(4), D
         => CoreAPB3_0_APBmslave0_PADDR(1), Y => \un5_penable_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_1_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    \fsmsync_ns_i_1[6]\ : CFG4
      generic map(INIT => x"F7F4")

      port map(A => \SDAInt\, B => \fsmsync[1]_net_1\, C => 
        N_1002, D => N_997, Y => \fsmsync_ns_i_1[6]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => N_1449, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_1_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[16]_net_1\, 
        C => \fsmsta[20]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_2181, B => N_145, C => N_166, D => 
        fsmsta_8_20_379_i_0_o2_0, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_sm0, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[15]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[6]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_9_509_0_1, D => N_1717, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_126, B => N_80, C => un136_framesync, Y => 
        N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => un92_fsmsta, B => un105_ens1, C => 
        \serdat_i_m_1[7]\, D => bsd7_tmp_i_m_1, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \PCLKint\, B => \un151_framesync\, C => 
        \PCLKint_ff\, Y => \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \fsmmod_ns_0_a4_0[5]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => N_1044, 
        D => un115_fsmdet, Y => N_1059);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \fsmsync_ns_i_o3_0[6]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => un70_fsmsta, B => \fsmsync[5]_net_1\, C => 
        N_64, Y => N_995);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => N_145_2, Y => fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[4]_net_1\, C => N_1727_2, 
        D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmmod_ns_0_a4_0_4[3]_net_1\, B => 
        un115_fsmdet, C => \fsmmod[3]_net_1\, D => N_1034, Y => 
        \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \sersta_32_2[0]\, B => N_72_mux, C => N_127, 
        D => \sersta_32_3[0]\, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un135_ens1_4, B => un135_ens1_5, C => 
        \un1_fsmsta_1_i_0_o2_0\, D => un135_ens1_3, Y => 
        un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0031")

      port map(A => \fsmmod[6]_net_1\, B => \fsmmod[2]_net_1\, C
         => \adrcomp\, D => \fsmmod[0]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3[19]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => \SDAInt\, B => N_2178, C => N_2177, D => 
        N_191, Y => N_157);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \un3_penable_1\, B => \un105_ens1_1\, C => 
        N_138, Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    \fsmsync_ns_i_a3_1_0_a2_2[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[3]_net_1\, C
         => \fsmmod[1]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\);
    
    \fsmmod_ns_0_o3[0]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => N_1040, B => \starto_en\, C => N_64, Y => 
        N_1044);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_1_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \fsmsync_RNO[1]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => N_995, B => \fsmsync_ns_i_1[6]_net_1\, C => 
        \fsmsync[1]_net_1\, D => \fsmsync[2]_net_1\, Y => 
        N_976_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_1656, B => \fsmdet[1]_net_1\, Y => N_1727_2);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => un115_fsmdet, B => N_1059, C => 
        \fsmmod[1]_net_1\, D => un10_sclscl, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_1_INT[0]\, 
        C => \fsmsta[28]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \serCON_WRITE_PROC.sercon_8_0_2[3]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \COREI2C_0_1_INT[0]\, B => N_163, C => N_162, 
        D => N_160, Y => \sercon_8_0_2[3]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_1_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[3]\ : CFG4
      generic map(INIT => x"6F60")

      port map(A => CO2_0, B => \framesync[3]_net_1\, C => 
        framesync_7_e2, D => \framesync_7_m2[3]\, Y => 
        \framesync_7[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    PCLK_count1_1_sqmuxa_1 : CFG4
      generic map(INIT => x"8CCC")

      port map(A => bclke, B => PCLK_count2_ov_6_1, C => 
        \sercon[7]_net_1\, D => \PCLK_count1_ov_1_sqmuxa_0\, Y
         => \PCLK_count1_1_sqmuxa_1\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[5]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG4
      generic map(INIT => x"0307")

      port map(A => \fsmmod[0]_net_1\, B => \nedetect\, C => 
        \fsmmod[4]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \fsmmod_ns_i_0[2]_net_1\);
    
    \FSMMOD_COMB_PROC.un10_sclscl\ : CFG2
      generic map(INIT => x"8")

      port map(A => \pedetect\, B => \SCLSCL\, Y => un10_sclscl);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_1586_1, B => N_2177, C => \fsmsta[8]_net_1\, 
        D => N_172, Y => fsmsta_8_5_555_a3_2);
    
    \fsmmod_ns_i_o3_0_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_1_INT[0]\, B => \sercon[4]_net_1\, 
        Y => N_997);
    
    adrcomp_2_sqmuxa_i_a3_2_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, C => \framesync[0]_net_1\, D => 
        \nedetect\, Y => \adrcomp_2_sqmuxa_i_a3_2_0\);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_0);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_0 is

    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          COREI2C_0_1_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          un3_penable                                : in    std_logic;
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_1_SCL_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_1_SDA_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          un3_penable_1                              : out   std_logic;
          un105_ens1_3                               : in    std_logic;
          un105_ens1_1                               : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic;
          un5_penable_1                              : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          bclke                                      : in    std_logic;
          N_138                                      : in    std_logic
        );

end COREI2C_0;

architecture DEF_ARCH of COREI2C_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_0
    port( COREI2C_0_1_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0) := (others => 'U');
          seradr0apb                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_1_SCL_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_1_SDA_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          un3_penable_1                              : out   std_logic;
          un105_ens1_3                               : in    std_logic := 'U';
          un105_ens1_1                               : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic := 'U';
          un5_penable_1                              : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          bclke                                      : in    std_logic := 'U';
          N_138                                      : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_0
	Use entity work.COREI2CREAL_6_0(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_0
      port map(COREI2C_0_1_SDAO_i(0) => COREI2C_0_1_SDAO_i(0), 
        COREI2C_0_1_SCLO_i(0) => COREI2C_0_1_SCLO_i(0), 
        COREI2C_0_1_INT(0) => COREI2C_0_1_INT(0), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, N_1221 => N_1221, N_1217 => 
        N_1217, N_1218 => N_1218, N_1220 => N_1220, N_1219 => 
        N_1219, BIBUF_COREI2C_0_1_SCL_IO_Y => 
        BIBUF_COREI2C_0_1_SCL_IO_Y, BIBUF_COREI2C_0_1_SDA_IO_Y
         => BIBUF_COREI2C_0_1_SDA_IO_Y, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, un3_penable_1 => 
        un3_penable_1, un105_ens1_3 => un105_ens1_3, un105_ens1_1
         => un105_ens1_1, CONFIG_rega20_2 => CONFIG_rega20_2, 
        un5_penable_1 => un5_penable_1, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, bclke => bclke, N_138 => 
        N_138);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_4 is

    port( COREI2C_0_5_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          seradr0apb                   : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          N_1218                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_5_SCL_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_5_SDA_IO_Y   : in    std_logic;
          bclke                        : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un105_ens1_0                 : in    std_logic;
          un105_ens1_3                 : in    std_logic;
          un3_penable_1                : in    std_logic;
          N_43                         : in    std_logic;
          un5_penable_0                : in    std_logic
        );

end COREI2CREAL_6_4;

architecture DEF_ARCH of COREI2CREAL_6_4 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_5_SDAO[0]\, \COREI2C_0_5_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_5_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        un1_serdat_2_sqmuxa_4, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, fsmsta_8_3_601, \fsmsta[9]_net_1\, 
        N_2172_i_0, \fsmsta[8]_net_1\, N_1665, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, fsmsta_8_13_406, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, fsmsta_8_28_307_0, \ack\, ack_7, 
        SDAO_int_7_0_275_0, SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, 
        bsd7_tmp_6, \bsd7\, bsd7_9_iv_i_0, \adrcomp\, N_2176, 
        adrcomp_2_sqmuxa_i_0_4, \PCLKint\, PCLKint_3, 
        un1_pclkint4_i_0, \ack_bit\, \ack_bit_1_sqmuxa\, 
        \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_4, un1_rtn_3_4, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, 
        \un1_PCLK_count1_0_sqmuxa_2\, 
        \un1_PCLK_count1_0_sqmuxa_3\, \PCLK_count1_ov_1_sqmuxa\, 
        PCLK_count2_ov_6_1, \un1_counter_rst_3\, N_997, 
        un70_fsmsta, N_1046, \fsmsta_cnst[0]\, N_1622_2, 
        \adrcomp_2_sqmuxa_i_o2_1_3\, N_66, N_84, N_1586_1, N_2181, 
        un105_ens1, \un1_serdat_2_sqmuxa_1_0\, un57_fsmsta, 
        \un1_serdat40\, N_2177, N_2173_i_1, N_133, un1_fsmmod, 
        N_36_i_1, un136_framesync, N_2196, N_2186, 
        \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, 
        \un1_pclk_count1_ov_1_1\, \un1_pclk_count1_ov_1\, N_23, 
        \sersta_32_1[2]\, \sersta_32_7[2]\, un135_ens1_2, 
        \un1_PCLK_count1_0_sqmuxa_0_1_0\, 
        \un1_PCLK_count1_0_sqmuxa_0\, \PRDATA_3_1_1[4]\, 
        \PRDATA_3_1_1[3]\, \PRDATA_3_1_1[7]\, \PRDATA_3_1_1[5]\, 
        \PRDATA_3_1_1[6]\, \fsmsta_8_ns_1[29]\, 
        \fsmsta_8_ns_1[28]\, \fsmsta_8_ns_1[16]\, un133_framesync, 
        un13_adrcompen, \fsmsta_8_ns_1[18]\, 
        \framesync_7_enl_bm_1[3]\, framesync_7_e2, 
        \framesync_7_enl_am_1[3]\, CO0, N_2179, N_1652, N_161_2, 
        fsmsta_8_5_555_a3_0_2, fsmsta_8_5_555_a3_2, 
        PCLK_count2_ov_6_0_a2_1_0, un111_fsmdet_0, 
        \sersta_32_i_a2_5[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, N_629, un139_ens1_0, 
        \adrcomp_2_sqmuxa_i_o2_1_1\, N_127, N_64, N_2178, N_1035, 
        N_67, N_153_1, N_26, un26_adrcompen_0, un10_sclscl, 
        N_1002_3, \un151_framesync\, N_1196, N_1197, N_1198, 
        SDAO_int_7_0_275_1, \adrcomp_2_sqmuxa_i_a3_3\, 
        SDAO_int_7_0_275_a5_0, un141_ens1_2, 
        \SDAO_int_1_sqmuxa_3\, \adrcomp_2_sqmuxa_i_a2_1_2\, 
        \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_10_476_i_a6_1, 
        \fsmmod_ns_i_a4_1_0[2]_net_1\, \sersta_32_4[0]\, 
        \sersta_32_3[0]\, \sersta_32_5[1]\, \sersta_32_4[1]\, 
        fsmsta_8_20_379_i_0_a3_5, fsmsta_8_20_379_i_0_a3_4, 
        \sersta_32_i_a2_7[4]\, \sersta_32_i_a2_6[4]\, 
        \sersta_32_4[2]\, un135_ens1_5, un135_ens1_3, 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0, 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0, un25_fsmsta_2, 
        \sersta_32_i_a2_8[3]\, \sersta_32_i_a2_7[3]\, 
        un13_adrcompen_4, m7_5, m7_4, N_1064, un33_fsmsta, 
        framesync_7_sm0, PCLK_count2_ov_6_0_a2_1_4_tz, N_1034, 
        N_2182, N_76, N_95, un16_fsmmod, CO2, 
        \un1_pclk_count1_ov\, CO1, N_1717, 
        \adrcomp_2_sqmuxa_i_a3_4\, \fsmmod_ns_i_0[2]_net_1\, 
        fsmsta_8_10_476_i_0, \SDAO_int_1_sqmuxa_4\, 
        \adrcomp_2_sqmuxa_i_a2_1_4\, PCLK_count2_ov_6_0_a2_1_3, 
        \sercon_8_2[4]\, fsmsta_8_3_601_a4_0_2, 
        \sersta_32_i_a2_9[4]\, un135_ens1_7_0, 
        fsmsta_8_9_509_a4_0_1, \sersta_32_i_a2_10[3]\, 
        un25_fsmsta, N_104, N_1044, un25_framesync, 
        un19_framesync, N_1002, N_2192, \fsmsta_8_0_a2_1[7]\, 
        N_1656, N_1041, N_130, N_995, N_191, N_2193, un74_ens1, 
        N_63, \un1_pclk_count191\, un23_pclk_count1, N_2171, 
        \un1_fsmsta_6\, N_1659_2, N_124, N_120, 
        fsmsta_8_28_307_a3_0_1, \SDAO_int_1_sqmuxa_7\, 
        \fsmsync_ns_i_1[6]_net_1\, \adrcomp_2_sqmuxa_i_a2_1_5\, 
        N_163, un135_ens1, N_162, N_165, \fsmsta_nxt_9_m[22]\, 
        \fsmsta_nxt_9_m[27]\, N_157, \framesync_1_sqmuxa\, N_1054, 
        un115_fsmdet, \fsmsta_nxt_9_m[26]\, \fsmsta_nxt_9_m[21]\, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, N_2188, N_160, N_1060, 
        N_1624, N_1657_2, N_70, \PCLK_count1_0_sqmuxa_3\, N_126, 
        \fsmsta_8_i_0[25]\, fsmsta_8_4_577_i_0, N_1729, N_1659, 
        N_82, N_80, bsd7_i_m_0, bsd7_tmp_i_m_2, 
        \fsmmod_ns_0_0[0]_net_1\, fsmsta_8_20_379_i_0_o2_0, 
        \un1_PCLK_count1_0_sqmuxa_1\, fsmsta_8_23_351_i_0_1, 
        \fsmsync_ns_0_0_1[0]_net_1\, 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\, N_1727, N_145, N_166, 
        N_1465, N_1657, \fsmsync_ns_i_0_1_tz[3]_net_1\, N_2198, 
        N_86, un1_fsmsta_10_i_0, N_2199, \PWDATA_i_m_1[7]\, 
        \sercon_8_0_2[3]\, N_1059, N_1486, N_1051, 
        \serdat_2_sqmuxa_0\, CO1_0, N_161, un134_fsmsta, 
        \serdat_0_sqmuxa\, \framesync_7_m2[3]\, N_2187, N_1466, 
        bsd7_tmp_6_sn_N_10_mux, bsd7_tmp_6_m1, bsd7_tmp_6_sm0, 
        CO0_0, bsd7_9_iv_1, CO1_1, bsd7_i_m, 
        \un1_serdat_2_sqmuxa_1\ : std_logic;

begin 

    COREI2C_0_5_INT(0) <= \COREI2C_0_5_INT[0]\;

    un151_framesync_RNIAL6C1 : CFG3
      generic map(INIT => x"DC")

      port map(A => \un151_framesync\, B => N_2177, C => N_191, Y
         => un1_fsmsta_10_i_0);
    
    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    adrcomp_2_sqmuxa_i_0_0 : CFG4
      generic map(INIT => x"0015")

      port map(A => un16_fsmmod, B => N_2192, C => 
        \COREI2C_0_5_INT[0]\, D => N_1586_1, Y => N_2176);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_153_1, 
        Y => N_2171);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_191, B => \un1_fsmsta_6\, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => N_166);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \framesync_7_enl_bm_1[3]\, B => 
        framesync_7_e2, C => \framesync_7_enl_am_1[3]\, Y => 
        \framesync_7[3]\);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[10]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[1]_net_1\, B => seradr0apb(2), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_0, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_4, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \bsd7\, Y => bsd7_i_m_0);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_1656, B => \fsmdet[1]_net_1\, Y => N_1657_2);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[14]_net_1\, 
        C => un25_fsmsta_2, D => N_2178, Y => un25_fsmsta);
    
    \fsmmod_ns_0_a4_0[1]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => N_1044, 
        D => un115_fsmdet, Y => N_1051);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \fsmsta[25]_net_1\, B => N_23, C => 
        \sersta_32_1[2]\, D => \sersta_32_7[2]\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, B => 
        \sercon[4]_net_1\, C => N_1041, D => N_1035, Y => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    un7_fsmsta_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[22]_net_1\, 
        Y => N_2178);
    
    \fsmmod_ns_0[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un115_fsmdet, B => \fsmmod_ns_0_0[0]_net_1\, 
        C => N_1064, Y => \fsmmod_ns[0]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    \fsmmod_ns_0_0[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => N_1044, D => un10_sclscl, Y => 
        \fsmmod_ns_0_0[0]_net_1\);
    
    PCLKint_ff_RNIODJV : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_1\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_2181, B => \adrcompen\, C => N_26, Y => 
        fsmsta_8_28_307_a3_0_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => un1_fsmmod, B => SDAO_int_7_0_275_1, C => 
        SDAO_int_7_0_275_a5_0, D => N_1466, Y => 
        SDAO_int_7_0_275_0);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \fsmsta_cnst[0]\, B => N_1657_2, C => 
        \fsmsta[4]_net_1\, D => \fsmdet[3]_net_1\, Y => N_1657);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CEFF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \un1_pclk_count1_ov_1_1\, D => 
        \sercon[7]_net_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => un139_ens1_0, Y => 
        framesync_7_sm0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"003A")

      port map(A => \ack\, B => N_172, C => N_2177, D => 
        fsmsta_8_4_577_i_0, Y => N_2172_i_0);
    
    un1_PCLK_count1_0_sqmuxa_0 : CFG4
      generic map(INIT => x"0031")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \sercon[1]_net_1\, C => \un1_PCLK_count1_0_sqmuxa_0_1_0\, 
        D => \sercon[7]_net_1\, Y => \un1_PCLK_count1_0_sqmuxa_0\);
    
    \fsmsta_RNO[25]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => N_172, B => N_2177, C => \fsmsta_8_i_0[25]\, 
        D => un136_framesync, Y => N_2175_i_0);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync[2]_net_1\, D => \framesync[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \fsmsta[17]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_2[3]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \sercon[6]_net_1\, B => \adrcomp\, C => 
        N_1586_1, D => un74_ens1, Y => N_163);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1652, Y => N_1656);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_RNIQ5T41\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \nedetect\, B => \COREI2C_0_5_INT[0]\, C => 
        un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sn_N_10_mux);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_5_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        N_161_2, Y => N_161);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \un1_PCLK_count1_1.CO1\ : CFG4
      generic map(INIT => x"8880")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_PCLK_count1_0_sqmuxa_2\, 
        D => \un1_PCLK_count1_0_sqmuxa_3\, Y => CO1_1);
    
    \serdat_RNIFRN01[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_5_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_66, B => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"FE0E")

      port map(A => \sercon_8_0_2[3]\, B => N_161, C => 
        un5_penable, D => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \sercon_9[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[18]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    SCLO_int_RNICG37 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_5_SCLO[0]\, Y => 
        COREI2C_0_5_SCLO_i(0));
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_4);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6s2\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_5_INT[0]\, 
        C => un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sm0);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmsta_cnst[0]\, D => \sercon[6]_net_1\, Y => 
        \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_5_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \un1_PCLK_count1_1.CO0\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \un1_PCLK_count1_0_sqmuxa_2\, C => 
        \un1_PCLK_count1_0_sqmuxa_3\, Y => CO0_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"D555")

      port map(A => N_2176, B => N_2187, C => N_95, D => 
        \adrcomp_2_sqmuxa_i_a3_4\, Y => adrcomp_2_sqmuxa_i_0_4);
    
    \un2_framesync_1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync_1_sqmuxa\, C => \framesync[1]_net_1\, Y => 
        CO1_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_629, B => \fsmmod[2]_net_1\, Y => 
        SDAO_int_7_0_275_a5_0);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \COREI2C_0_5_SDAO[0]\, B => N_2177, C => 
        fsmsta_8_23_351_i_0_1, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \fsmsync_ns_0_a3_2_2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[4]_net_1\, Y
         => N_1002_3);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0045")

      port map(A => bsd7_9_iv_1, B => \serdat[7]_net_1\, C => 
        bsd7_tmp_6_sn_N_10_mux, D => bsd7_i_m, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[0]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    \sersta_RNIAMG52[4]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        \sercon[7]_net_1\, Y => N_1221);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    un1_fsmsta_nxt_0_sqmuxa_i_a3_1 : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, Y
         => N_153_1);
    
    \serCON_WRITE_PROC.sercon_8_0_a3[3]\ : CFG4
      generic map(INIT => x"CC08")

      port map(A => \fsmdet[3]_net_1\, B => \sercon[6]_net_1\, C
         => N_629, D => N_1064, Y => N_160);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_11_454_i_a6_2_0_0_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, Y => 
        N_2182);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_0, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[12]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2177, B => N_2178, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, Y
         => N_629);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    framesync_1_sqmuxa : CFG3
      generic map(INIT => x"20")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, Y
         => \framesync_1_sqmuxa\);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_5_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    un1_fsmsta_1_i_0_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[12]_net_1\, 
        C => \fsmsta[16]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => fsmsta_8_28_307_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    \serdat_RNIC6Q81[7]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(7), B => \serdat[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    un1_fsmsta_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[14]_net_1\, 
        C => \fsmsta[18]_net_1\, Y => N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[0]\ : CFG4
      generic map(INIT => x"6F60")

      port map(A => \framesync_1_sqmuxa\, B => 
        \framesync[0]_net_1\, C => framesync_7_e2, D => 
        \framesync_7_m2[3]\, Y => \framesync_7[0]\);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    \sersta_RNIU9G52[1]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[4]\, C => \sersta[1]_net_1\, D => 
        seradr0apb(4), Y => N_1218);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => fsmsta_8_3_601, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[26]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_18_s5_1_0, Y => 
        \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \CLK_COUNTER1_PROC.un1_bclke_1.CO2\ : CFG3
      generic map(INIT => x"01")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[21]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_RNIQK8M1[5]\ : CFG4
      generic map(INIT => x"FEF0")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmsta_cnst[0]\, D => \fsmdet[3]_net_1\, Y => 
        N_1622_2);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    serdat_2_sqmuxa_0 : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_5_INT[0]\, B => un57_fsmsta, C => 
        \fsmdet[3]_net_1\, Y => \serdat_2_sqmuxa_0\);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \COREI2C_0_5_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \ack\, B => N_2177, C => N_133, D => 
        fsmsta_8_28_307_a3_0_1, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \COREI2C_0_5_INT[0]\, D => \sersta_32_i_a2_7[3]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"0002")

      port map(A => PCLK_count2_ov_6_1, B => 
        \PCLK_count1_ov_1_sqmuxa\, C => 
        \un1_PCLK_count1_0_sqmuxa_3\, D => 
        \un1_PCLK_count1_0_sqmuxa_2\, Y => \PCLK_count1_1_sqmuxa\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[6]_net_1\, C
         => \fsmmod[1]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_5_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \un1_counter_rst_3\, D => 
        CO0_0, Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[16]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_1[3]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        N_2177, D => N_2179, Y => N_162);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[14]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmmod_ns_i_o3_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_5_INT[0]\, B => \sercon[5]_net_1\, 
        Y => N_1035);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"00D0")

      port map(A => N_2186, B => N_2177, C => N_82, D => 
        un136_framesync, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \sersta_RNIQ5G52[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"88A8")

      port map(A => \SCLInt\, B => \fsmdet[3]_net_1\, C => 
        \fsmdet[2]_net_1\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \sersta_32_4[1]\, B => m7_4, C => 
        \sersta_32_5[1]\, D => m7_5, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNI3GU11 : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        un136_framesync, C => \pedetect\, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[27]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_24_s4_1_0, Y => 
        \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[3]\ : CFG4
      generic map(INIT => x"7F80")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, C => CO0, D => \framesync[3]_net_1\, 
        Y => \framesync_7_enl_bm_1[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG3
      generic map(INIT => x"32")

      port map(A => fsmsta_8_5_555_a3_0_2, B => N_2181, C => 
        fsmsta_8_5_555_a3_2, Y => N_1665);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_5_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_5_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"54F0")

      port map(A => \ack\, B => seradr0apb(0), C => 
        \adrcomp_2_sqmuxa_i_a2_1_5\, D => un13_adrcompen, Y => 
        N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => fsmsta_8_13_406);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_5_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7[0]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_m2[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => fsmsta_8_28_307_0);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \fsmsta_RNO[19]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_2199, B => un136_framesync, C => N_157, Y
         => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => fsmsta_8_13_406, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_PCLK_count1_0_sqmuxa_0_1_0 : CFG4
      generic map(INIT => x"577F")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count1[1]_net_1\, D => 
        \PCLK_count1[0]_net_1\, Y => 
        \un1_PCLK_count1_0_sqmuxa_0_1_0\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_1041, B => N_1035, C => 
        \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => N_1054);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_0\ : CFG4
      generic map(INIT => x"CFEE")

      port map(A => N_2182, B => N_2181, C => \fsmsta[9]_net_1\, 
        D => N_2177, Y => fsmsta_8_4_577_i_0);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    \sercon_RNIJVN01[5]\ : CFG4
      generic map(INIT => x"05F3")

      port map(A => \serdat[5]_net_1\, B => \sercon[5]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[5]\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFDC")

      port map(A => N_2177, B => un16_fsmmod, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \fsmsta[11]_net_1\, B => N_2177, C => N_120, 
        Y => N_2198);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_5_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO0, B => framesync_7_e2, C => 
        \framesync[1]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[1]\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => un16_fsmmod, B => \sercon_8_2[4]\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), D => un5_penable, Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_76, Y => N_55_i_0);
    
    un1_PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"CCEF")

      port map(A => CO2, B => \un1_PCLK_count1_0_sqmuxa_1\, C => 
        \PCLK_count1[3]_net_1\, D => \sercon[7]_net_1\, Y => 
        \un1_PCLK_count1_0_sqmuxa_3\);
    
    \FSMSTA_SYNC_PROC.un133_framesync\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \pedetect\, B => \fsmsta[23]_net_1\, C => 
        un1_fsmmod, D => N_2177, Y => un133_framesync);
    
    \serSTA_WRITE_PROC.sersta_32_1[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[24]_net_1\, B => \fsmsta[16]_net_1\, 
        C => \fsmsta[15]_net_1\, D => un135_ens1_2, Y => 
        \sersta_32_1[2]\);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un133_framesync, B => N_2181, Y => 
        un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0056")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \un1_PCLK_count1_0_sqmuxa_2\, C => 
        \un1_PCLK_count1_0_sqmuxa_3\, D => \un1_counter_rst_3\, Y
         => \PCLK_count1_10[0]\);
    
    \serSTA_WRITE_PROC.sersta_32_4[0]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => \COREI2C_0_5_INT[0]\, B => N_127, C => 
        \fsmsta[9]_net_1\, Y => \sersta_32_4[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO\ : CFG4
      generic map(INIT => x"C010")

      port map(A => \nedetect\, B => \COREI2C_0_5_INT[0]\, C => 
        bsd7_i_m_0, D => un105_ens1, Y => bsd7_i_m);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    un1_PCLK_count1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"CECC")

      port map(A => bclke, B => \PCLK_count1_0_sqmuxa_3\, C => 
        \PCLK_count1[3]_net_1\, D => CO2, Y => 
        \un1_PCLK_count1_0_sqmuxa_1\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG3
      generic map(INIT => x"37")

      port map(A => N_67, B => \fsmsync[4]_net_1\, C => N_66, Y
         => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    \un2_framesync_1_1.CO0\ : CFG3
      generic map(INIT => x"08")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        un70_fsmsta, Y => CO0);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_0_2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \adrcomp\, B => \framesync[0]_net_1\, C => 
        \framesync[3]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        fsmsta_8_3_601_a4_0_2);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"F7F5")

      port map(A => N_2178, B => \fsmsta[20]_net_1\, C => N_2188, 
        D => N_2177, Y => fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => \fsmmod[2]_net_1\, B => N_1064, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un5_penable_0, B => un105_ens1_3, C => 
        un3_penable_1, D => N_43, Y => un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"2220")

      port map(A => PCLK_count2_ov_6_0_a2_1_3, B => un16_fsmmod, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    SDAO_int_RNI2V2A : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_5_SDAO[0]\, Y => 
        COREI2C_0_5_SDAO_i(0));
    
    un1_counter_rst_3 : CFG4
      generic map(INIT => x"01FF")

      port map(A => \un1_PCLK_count1_0_sqmuxa_2\, B => 
        \un1_PCLK_count1_0_sqmuxa_3\, C => 
        \PCLK_count1_ov_1_sqmuxa\, D => PCLK_count2_ov_6_1, Y => 
        \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_5_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"CACC")

      port map(A => \COREI2C_0_5_SDAO[0]\, B => 
        \fsmsta[13]_net_1\, C => N_2177, D => N_2196, Y => N_82);
    
    \fsmsta_RNO[12]\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_124, B => N_2188, C => N_2186, Y => 
        N_1774_i_0);
    
    PCLK_count1_ov_1_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \sercon[7]_net_1\, B => bclke, C => 
        \sercon[1]_net_1\, D => \sercon[0]_net_1\, Y => 
        \PCLK_count1_ov_1_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_5_SDAO[0]\, Y => 
        N_172);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_m1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        \serdat_0_sqmuxa\, Y => bsd7_tmp_6_m1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_4, B => N_153_1, C => 
        N_2177, D => fsmsta_8_20_379_i_0_a3_5, Y => N_145);
    
    adrcomp : SLE
      port map(D => N_2176, CLK => FAB_CCC_GL0, EN => 
        adrcomp_2_sqmuxa_i_0_4, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[27]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_4);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \fsmdet[3]_net_1\, B => N_629, C => 
        \fsmdet[1]_net_1\, Y => N_1717);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_5\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => un135_ens1_2, Y => un135_ens1_5);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[7]_net_1\, C
         => \fsmsta[11]_net_1\, D => \fsmsta[9]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => \fsmsta[16]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        un25_fsmsta_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \PCLKint\, B => \PCLKint_ff\, C => N_1586_1, 
        D => \fsmmod[2]_net_1\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG3
      generic map(INIT => x"BF")

      port map(A => N_997, B => un70_fsmsta, C => 
        \fsmmod[4]_net_1\, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[26]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_0_1\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \adrcomp\, B => \framesync[0]_net_1\, C => 
        \framesync[3]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        fsmsta_8_9_509_a4_0_1);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => N_1665, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    un1_PCLK_count1_0_sqmuxa_2 : CFG4
      generic map(INIT => x"CCCE")

      port map(A => un23_pclk_count1, B => 
        \un1_PCLK_count1_0_sqmuxa_0\, C => \sercon[0]_net_1\, D
         => \sercon[7]_net_1\, Y => \un1_PCLK_count1_0_sqmuxa_2\);
    
    \sersta_RNI2EG52[2]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        seradr0apb(5), Y => N_1219);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \fsmsync[5]_net_1\, B => N_64, C => 
        \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \fsmmod[5]_net_1\, B => \nedetect\, C => 
        un115_fsmdet, D => N_1051, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_5_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => un135_ens1_2, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG4
      generic map(INIT => x"2220")

      port map(A => N_2198, B => N_2188, C => \fsmsta[11]_net_1\, 
        D => N_2186, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_3\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[8]_net_1\, B => \fsmsta[16]_net_1\, C
         => \fsmsta[20]_net_1\, D => \fsmsta[2]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[22]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[22]\, Y => 
        \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_4, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG3
      generic map(INIT => x"06")

      port map(A => \PCLK_count1[1]_net_1\, B => CO0_0, C => 
        \un1_counter_rst_3\, Y => \PCLK_count1_10[1]\);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_64, D => N_1002_3, Y => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \bsd7_tmp\, B => \SCLInt\, C => 
        \COREI2C_0_5_INT[0]\, D => un57_fsmsta, Y => 
        bsd7_tmp_i_m_2);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"F0F8")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat_2_sqmuxa_1_0\, Y => 
        un1_serdat_2_sqmuxa_4);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \indelay[1]_net_1\, B => \indelay[3]_net_1\, 
        Y => N_66);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \fsmsta_cnst[0]\, B => N_1657_2, C => 
        \fsmsta[10]_net_1\, D => \fsmdet[3]_net_1\, Y => N_1727);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1002, B => \COREI2C_0_5_INT[0]\, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_5_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FF7F")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_66, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_5_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"0C08")

      port map(A => \serdat_2_sqmuxa_0\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_7\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, D => un135_ens1_5, Y => 
        un135_ens1_7_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_26_328_a3_0_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => \fsmsta[23]_net_1\, B => \adrcomp\, Y => N_26);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1717, B => fsmsta_8_3_601_a4_0_2, C => 
        N_1729, D => N_1727, Y => fsmsta_8_3_601);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_172, B => N_2182, C => N_2193, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_1002_3, B => 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[2]_net_1\, Y => N_1002);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[27]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => \serdat[3]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[7]_net_1\, C
         => \fsmsta[11]_net_1\, D => \fsmsta[23]_net_1\, Y => 
        m7_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[26]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_1\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \adrcomp\, B => \framesync[3]_net_1\, C => 
        N_1652, D => N_1659_2, Y => N_1729);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ack\, B => \adrcompen\, C => N_2177, D => 
        N_26, Y => fsmsta_8_5_555_a3_0_2);
    
    \sersta_RNI6IG52[3]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        \sercon[6]_net_1\, Y => N_1220);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_5_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3340")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1586_1, Y => N_1624);
    
    adrcomp_2_sqmuxa_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[23]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => N_95);
    
    serdat_0_sqmuxa : CFG3
      generic map(INIT => x"08")

      port map(A => \COREI2C_0_5_INT[0]\, B => un57_fsmsta, C => 
        \fsmdet[3]_net_1\, Y => \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        \COREI2C_0_5_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_1046, B => \fsmmod_ns_i_0[2]_net_1\, C => 
        N_1054, D => un115_fsmdet, Y => N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[23]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_5);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_o3\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2181, B => N_1656, Y => N_2188);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_5_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \serdat_RNIHTN01[4]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[4]_net_1\, B => \sercon[4]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[4]\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    \fsmsync_ns_i_1[6]\ : CFG4
      generic map(INIT => x"F7F4")

      port map(A => \SDAInt\, B => \fsmsync[1]_net_1\, C => 
        N_1002, D => N_997, Y => \fsmsync_ns_i_1[6]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(4), B => seradr0apb(3), C => 
        \serdat[3]_net_1\, D => \serdat[2]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => SDAO_int_7_0_275_0, CLK => FAB_CCC_GL0, EN
         => SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \COREI2C_0_5_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[19]_net_1\, 
        C => \fsmsta[16]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_2181, B => N_145, C => 
        fsmsta_8_20_379_i_0_o2_0, D => N_166, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_sm0, Y => framesync_7_e2);
    
    \serdat_RNIA4Q81[6]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(6), B => \serdat[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[6]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[15]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[2]_net_1\, B => \serdat[1]_net_1\, C
         => \serdat[0]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    \fsmsync_ns_i_a3_1_0_a2_1[2]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, Y
         => \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \fsmsta_RNO[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_126, B => N_80, C => un136_framesync, Y => 
        N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"FBF8")

      port map(A => \PWDATA_i_m_1[7]\, B => un105_ens1, C => 
        \fsmdet[3]_net_1\, D => bsd7_tmp_i_m_2, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \PCLKint\, B => \un151_framesync\, C => 
        \PCLKint_ff\, Y => \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \fsmmod_ns_0_a4_0[5]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \fsmmod[6]_net_1\, B => \SDAInt\, C => N_1044, 
        D => un115_fsmdet, Y => N_1059);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \fsmsync_ns_i_o3_0[6]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => un70_fsmsta, B => \fsmsync[5]_net_1\, C => 
        N_64, Y => N_995);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_1\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \adrcomp\, B => \framesync[3]_net_1\, C => 
        N_1652, D => N_1659_2, Y => N_1659);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[0]_net_1\, B => seradr0apb(1), Y => 
        un26_adrcompen_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => N_1659, B => N_1657, C => N_1717, D => 
        fsmsta_8_9_509_a4_0_1, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"5444")

      port map(A => un115_fsmdet, B => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, C => \fsmmod[3]_net_1\, D
         => N_1034, Y => \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FDFF")

      port map(A => m7_4, B => \sersta_32_3[0]\, C => 
        \sersta_32_4[0]\, D => m7_5, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        C => un135_ens1_7_0, D => un135_ens1_3, Y => un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_4, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0301")

      port map(A => \fsmmod[6]_net_1\, B => \fsmmod[2]_net_1\, C
         => \fsmmod[0]_net_1\, D => \adrcomp\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_1_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_1717, B => \fsmsta_cnst[0]\, Y => N_1659_2);
    
    un1_serdat_2_sqmuxa_1_0 : CFG4
      generic map(INIT => x"00EF")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_5_INT[0]\, 
        C => un57_fsmsta, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1_0\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => \bsd7_tmp\, B => bsd7_tmp_6_m1, C => 
        bsd7_tmp_6_sm0, D => bsd7_tmp_6_sn_N_10_mux, Y => 
        bsd7_tmp_6);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3[19]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => \SDAInt\, B => N_2178, C => N_2177, D => 
        N_191, Y => N_157);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un105_ens1_0, B => un105_ens1_3, C => 
        un3_penable_1, D => N_43, Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    \fsmmod_ns_0_o3[0]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \sercon[4]_net_1\, B => \starto_en\, C => 
        N_1035, D => N_64, Y => N_1044);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_5_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \fsmsync_RNO[1]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => N_995, B => \fsmsync_ns_i_1[6]_net_1\, C => 
        \fsmsync[1]_net_1\, D => \fsmsync[2]_net_1\, Y => 
        N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => un115_fsmdet, B => N_1059, C => 
        \fsmmod[1]_net_1\, D => un10_sclscl, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_5_INT[0]\, 
        C => \fsmsta[28]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \serCON_WRITE_PROC.sercon_8_0_2[3]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \COREI2C_0_5_INT[0]\, B => N_163, C => N_162, 
        D => N_160, Y => \sercon_8_0_2[3]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_5_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[3]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_enl_am_1[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[5]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG4
      generic map(INIT => x"0307")

      port map(A => \fsmmod[0]_net_1\, B => \nedetect\, C => 
        \fsmmod[4]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \fsmmod_ns_i_0[2]_net_1\);
    
    \FSMMOD_COMB_PROC.un10_sclscl\ : CFG2
      generic map(INIT => x"8")

      port map(A => \pedetect\, B => \SCLSCL\, Y => un10_sclscl);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_1586_1, B => N_2177, C => \fsmsta[8]_net_1\, 
        D => N_172, Y => fsmsta_8_5_555_a3_2);
    
    \fsmmod_ns_i_o3_0_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_5_INT[0]\, B => \sercon[4]_net_1\, 
        Y => N_997);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0_RNIN5VJ\ : CFG2
      generic map(INIT => x"1")

      port map(A => un57_fsmsta_1_0, B => N_2178, Y => N_191);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1_1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_4);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    
    \CLK_COUNTER1_PROC.un23_pclk_count1_1.CO3\ : CFG4
      generic map(INIT => x"3777")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => un23_pclk_count1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_4 is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          COREI2C_0_5_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          un3_penable                  : in    std_logic;
          N_1218                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_5_SCL_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_5_SDA_IO_Y   : in    std_logic;
          bclke                        : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un105_ens1_0                 : in    std_logic;
          un105_ens1_3                 : in    std_logic;
          un3_penable_1                : in    std_logic;
          N_43                         : in    std_logic;
          un5_penable_0                : in    std_logic
        );

end COREI2C_4;

architecture DEF_ARCH of COREI2C_4 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_4
    port( COREI2C_0_5_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          seradr0apb                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          N_1218                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_5_SCL_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_5_SDA_IO_Y   : in    std_logic := 'U';
          bclke                        : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un105_ens1_0                 : in    std_logic := 'U';
          un105_ens1_3                 : in    std_logic := 'U';
          un3_penable_1                : in    std_logic := 'U';
          N_43                         : in    std_logic := 'U';
          un5_penable_0                : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_4
	Use entity work.COREI2CREAL_6_4(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_4
      port map(COREI2C_0_5_SDAO_i(0) => COREI2C_0_5_SDAO_i(0), 
        COREI2C_0_5_SCLO_i(0) => COREI2C_0_5_SCLO_i(0), 
        COREI2C_0_5_INT(0) => COREI2C_0_5_INT(0), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, N_1218 => N_1218, N_1217 => 
        N_1217, N_1221 => N_1221, N_1219 => N_1219, N_1220 => 
        N_1220, BIBUF_COREI2C_0_5_SCL_IO_Y => 
        BIBUF_COREI2C_0_5_SCL_IO_Y, BIBUF_COREI2C_0_5_SDA_IO_Y
         => BIBUF_COREI2C_0_5_SDA_IO_Y, bclke => bclke, N_1214
         => N_1214, N_1215 => N_1215, N_1216 => N_1216, 
        un105_ens1_0 => un105_ens1_0, un105_ens1_3 => 
        un105_ens1_3, un3_penable_1 => un3_penable_1, N_43 => 
        N_43, un5_penable_0 => un5_penable_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity M2sExt_sb_CCC_0_FCCC is

    port( IO_0_Y       : in    std_logic_vector(0 to 0);
          FAB_CCC_GL0  : out   std_logic;
          FAB_CCC_LOCK : out   std_logic
        );

end M2sExt_sb_CCC_0_FCCC;

architecture DEF_ARCH of M2sExt_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => FAB_CCC_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FA0000045564000318C6318C1F18C61F00404040400403",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => IO_0_Y(0), CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        GND_net_1, RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_5 is

    port( COREI2C_0_6_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 2);
          seradr0apb                                 : in    std_logic_vector(7 downto 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          bclke                                      : in    std_logic;
          N_1218                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          BIBUF_COREI2C_0_6_SCL_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_6_SDA_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_8_0                                      : in    std_logic;
          un105_ens1_1                               : in    std_logic;
          un5_penable_1                              : in    std_logic
        );

end COREI2CREAL_6_5;

architecture DEF_ARCH of COREI2CREAL_6_5 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_6_SDAO[0]\, \COREI2C_0_6_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_6_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        un1_serdat_2_sqmuxa_5, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, N_1665, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, N_1470, \ack\, ack_7, N_1449, 
        SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, bsd7_tmp_6, \bsd7\, 
        bsd7_9_iv_i_0, \adrcomp\, N_2176, adrcomp_2_sqmuxa_i_0_5, 
        \PCLKint\, PCLKint_3, un1_pclkint4_i_0, \ack_bit\, 
        \ack_bit_1_sqmuxa\, \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_5, un1_rtn_3_5, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, 
        \PCLK_count1_ov_1_sqmuxa\, PCLK_count2_ov_6_1, 
        \PCLK_count1_1_sqmuxa_4\, \un1_counter_rst_3\, N_2177, 
        N_191, \un151_framesync\, un1_fsmsta_10_i_0, N_193, 
        N_1041, N_1043, N_997, un57_fsmsta, \un1_serdat40\, 
        \un1_serdat_2_sqmuxa_1_0\, \fsmsta_cnst[0]\, N_1622_2, 
        N_2182, ANC2, N_1586_1, N_2181, N_2173_i_1, N_133, 
        un1_fsmmod, N_36_i_1, un136_framesync, N_2196, N_2186, 
        \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, N_1717, N_1652, 
        fsmsta_8_9_509_0_1, fsmsta_8_9_509_0, fsmsta_8_3_601_0_1, 
        fsmsta_8_3_601_0, \un1_pclk_count1_ov_1_1\, 
        \un1_pclk_count1_ov_1\, \PCLK_count1_1_sqmuxa_1_0_1\, 
        \PCLK_count1_1_sqmuxa_1_0\, CO1, \PRDATA_3_1_1[4]\, 
        \PRDATA_3_1_1[7]\, \PRDATA_3_1_1[5]\, \PRDATA_3_1_1[3]\, 
        \PRDATA_3_1_1[6]\, un105_ens1, \fsmsta_8_ns_1[28]\, 
        \fsmsta_8_ns_1[29]\, \fsmsta_8_ns_1[16]\, un137_framesync, 
        un13_adrcompen, \fsmsta_8_ns_1[18]\, 
        \framesync_7_enl_bm_2[3]\, \framesync_7_enl_am_2[3]\, 
        framesync_7_e2, \framesync_7_enl_bm[0]\, 
        \framesync_7_enl_am[0]\, N_2171, \fsmsta_8_0_a2_1[7]\, 
        fsmsta_8_5_555_a3_0_2, fsmsta_8_5_555_a3_2, 
        PCLK_count2_ov_6_0_a2_1_1, un111_fsmdet_0, 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, 
        \adrcomp_2_sqmuxa_i_a3_1\, N_629, un139_ens1_0, 
        \adrcomp_2_sqmuxa_i_o2_1_1\, N_64, N_67, un135_ens1_2, 
        N_92, N_26, un135_ens1_7, un10_sclscl, CO1_0, un1_ens1, 
        un26_adrcompen_6, N_1002_3, N_1196, N_1197, N_1198, 
        un3_penable_0, \adrcomp_2_sqmuxa_i_a3_3\, un141_ens1_2, 
        \SDAO_int_1_sqmuxa_3\, \adrcomp_2_sqmuxa_i_a2_1_2\, 
        \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_10_476_i_a6_1, 
        \sersta_32_4[0]\, \sersta_32_3[0]\, \sersta_32_5[1]\, 
        \sersta_32_4[1]\, \fsmmod_ns_i_a4_1_0[2]_net_1\, 
        fsmsta_8_20_379_i_0_a3_4, fsmsta_8_20_379_i_0_a3_3_0, 
        \sersta_32_i_a2_8[4]\, \sersta_32_i_a2_7[4]\, 
        \sersta_32_i_a2_6[4]\, \sersta_32_i_a2_5[4]\, 
        \sersta_32_6[2]\, \sersta_32_5[2]\, \sersta_32_4[2]\, 
        \sersta_32_3[2]\, un135_ens1_5, un135_ens1_3, 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0, 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0, un25_fsmsta_1, 
        \sersta_32_i_a2_9[3]\, \sersta_32_i_a2_8[3]\, 
        \sersta_32_i_a2_7[3]\, \sersta_32_i_a2_6[3]\, 
        \adrcomp_2_sqmuxa_i_o2_1_2\, m7_4, m7_3, 
        \PCLK_count1_0_sqmuxa_4_1\, un13_adrcompen_4, N_1064, 
        framesync_7_e2_1, un33_fsmsta, 
        PCLK_count2_ov_6_0_a2_1_4_tz, un70_fsmsta, N_76, N_1040, 
        \un1_pclk_count1_ov\, CO1_1, N_1034, N_95, N_2179, 
        un16_fsmmod, \adrcomp_2_sqmuxa_i_a3_4\, 
        \fsmmod_ns_i_0[2]_net_1\, fsmsta_8_10_476_i_0, 
        \SDAO_int_1_sqmuxa_4\, \adrcomp_2_sqmuxa_i_a2_1_4\, 
        PCLK_count2_ov_6_0_a2_1_3, \fsmsta_8_i_a3_0[19]\, 
        \sercon_8_2[4]\, un135_ens1_7_0, N_104, un25_fsmsta, 
        un19_framesync, un25_framesync, N_2192, N_1002, N_995, 
        N_130, N_63, N_84, \un1_fsmsta_6\, un91_ens1, N_2193, 
        N_1656, un74_ens1, \un1_pclk_count191\, N_134, N_120, 
        N_124, fsmsta_8_28_307_a3_0_1, fsmsta_8_9_509_a4_0, 
        fsmsta_8_3_601_a4_0, \SDAO_int_1_sqmuxa_7\, 
        \fsmsync_ns_i_1[6]_net_1\, \adrcomp_2_sqmuxa_i_a2_1_5\, 
        fsmsta_8_20_379_i_0_a3_6, un135_ens1, 
        \fsmsta_nxt_9_m[26]\, \fsmsta_nxt_9_m[22]\, 
        \fsmsta_nxt_9_m[21]\, un115_fsmdet, N_165, N_1054, 
        \PCLK_count1_0_sqmuxa_1\, \fsmsta_nxt_9_m[27]\, N_163, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, N_1046, N_70, N_1624, 
        N_126, N_1048, \PCLK_count1_0_sqmuxa_2\, 
        \PCLK_count1_0_sqmuxa_3\, N_1060, \fsmsta_8_i_0[25]\, 
        fsmsta_8_4_577_i_0, N_80, N_82, bsd7_i_m_0, 
        bsd7_tmp_i_m_2, \PCLK_count1_1_sqmuxa_0\, 
        fsmsta_8_20_379_i_0_o2_0, \sercon_8_0_1[3]\, 
        \fsmsync_ns_0_0_1[0]_net_1\, fsmsta_8_23_351_i_0_1, 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\, N_1465, N_1058, N_1050, 
        \fsmsync_ns_i_0_1_tz[3]_net_1\, N_86, un92_fsmsta, CO0, 
        N_161_2, N_1059_1, N_2199, \PWDATA_i_m_1[7]\, 
        \sercon_8_0_2[3]\, fsmsta_8_2_647_i_0_0, N_91, N_1486, 
        \serdat_0_sqmuxa\, bsd7_tmp_6_m1, un134_fsmsta, N_2187, 
        CO1_2, N_161, N_1466, bsd7_tmp_6_sn_N_10_mux, CO0_0, 
        N_1467, bsd7_tmp_6_sm0, CO1_3, bsd7_9_iv_1, bsd7_i_m, 
        \un1_serdat_2_sqmuxa_1\ : std_logic;

begin 

    COREI2C_0_6_INT(0) <= \COREI2C_0_6_INT[0]\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG3
      generic map(INIT => x"40")

      port map(A => \framesync[3]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_a3_1\, C => \framesync[0]_net_1\, Y
         => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => N_2177, B => N_191, C => \un151_framesync\, Y
         => un1_fsmsta_10_i_0);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \sersta_32_i_a2_9[3]\, B => 
        \sersta_32_i_a2_7[3]\, C => \sersta_32_i_a2_6[3]\, D => 
        \sersta_32_i_a2_8[3]\, Y => N_99_i_0);
    
    adrcomp_2_sqmuxa_i_0_0 : CFG4
      generic map(INIT => x"0015")

      port map(A => un16_fsmmod, B => N_2192, C => 
        \COREI2C_0_6_INT[0]\, D => N_1586_1, Y => N_2176);
    
    \serdat_RNIA5801[5]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(5), B => \serdat[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmdet[1]_net_1\, B => \fsmsync[2]_net_1\, Y
         => PCLK_count2_ov_6_0_a2_1_1);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[0]_net_1\, B => seradr0apb(1), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG4
      generic map(INIT => x"CCCD")

      port map(A => \fsmsta[9]_net_1\, B => N_2177, C => 
        \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => N_2171);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_3\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[27]_net_1\, 
        C => \fsmsta[4]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_3);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \framesync_7_enl_bm_2[3]\, B => 
        \framesync_7_enl_am_2[3]\, C => framesync_7_e2, Y => 
        \framesync_7[3]\);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.CO1\ : CFG2
      generic map(INIT => x"7")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[0]_net_1\, Y => CO1_0);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[3]_net_1\, B => seradr0apb(4), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_6, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    \serSTA_WRITE_PROC.sersta_32_3[2]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \fsmsta[18]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => \fsmsta[26]_net_1\, Y => \sersta_32_3[2]\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_5, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \bsd7\, Y => bsd7_i_m_0);
    
    PCLK_count1_1_sqmuxa_4 : CFG4
      generic map(INIT => x"1000")

      port map(A => \PCLK_count1_0_sqmuxa_1\, B => 
        \PCLK_count1_0_sqmuxa_2\, C => \PCLK_count1_1_sqmuxa_1_0\, 
        D => \PCLK_count1_1_sqmuxa_0\, Y => 
        \PCLK_count1_1_sqmuxa_4\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[0]\ : CFG4
      generic map(INIT => x"C6CC")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        un70_fsmsta, D => N_2177, Y => \framesync_7_enl_bm[0]\);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_1);
    
    \fsmdet_RNIUR9P[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        C => un25_fsmsta_1, D => un135_ens1_7, Y => un25_fsmsta);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sersta_32_3[2]\, B => \sersta_32_6[2]\, C
         => \sersta_32_5[2]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1041, B => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, 
        C => N_1040, Y => \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    PCLK_count1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"0405")

      port map(A => \sercon[7]_net_1\, B => ANC2, C => 
        \sercon[0]_net_1\, D => \PCLK_count1[3]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_1\);
    
    \fsmmod_ns_0[0]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => N_1048, B => N_1043, C => \fsmmod[1]_net_1\, 
        D => un10_sclscl, Y => \fsmmod_ns[0]\);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \adrcomp_2_sqmuxa_i_o2_1_2\, D => 
        \adrcomp_2_sqmuxa_i_o2_1_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_1\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_2181, B => \adrcompen\, C => N_26, Y => 
        fsmsta_8_28_307_a3_0_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => \fsmmod[3]_net_1\, C
         => N_1467, D => un1_ens1, Y => N_1449);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \sercon[7]_net_1\, D => 
        \un1_pclk_count1_ov_1_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2\ : CFG4
      generic map(INIT => x"FF20")

      port map(A => \fsmsta[23]_net_1\, B => un1_fsmmod, C => 
        N_193, D => fsmsta_8_20_379_i_0_o2_0, Y => N_91);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"003A")

      port map(A => \ack\, B => N_172, C => N_2177, D => 
        fsmsta_8_4_577_i_0, Y => N_2172_i_0);
    
    \fsmsta_RNO[25]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => N_172, B => N_2177, C => \fsmsta_8_i_0[25]\, 
        D => un136_framesync, Y => N_2175_i_0);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_6\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), Y => 
        un26_adrcompen_6);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG3
      generic map(INIT => x"80")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \adrcomp_2_sqmuxa_i_a3_1\, Y => \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \fsmsta[17]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_2[3]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        N_1586_1, D => un74_ens1, Y => N_163);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1652, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG4
      generic map(INIT => x"008A")

      port map(A => \adrcomp\, B => \framesync[0]_net_1\, C => 
        \framesync[3]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        fsmsta_8_3_601_0_1);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \serdat_RNIH5T11[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_6_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_o2[3]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => N_1064, B => \fsmdet[3]_net_1\, C => N_629, Y
         => N_134);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_6_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        N_161_2, Y => N_161);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \un1_PCLK_count1_1.CO1\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \PCLK_count1_ov_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1[0]_net_1\, D => 
        \PCLK_count1[1]_net_1\, Y => CO1_3);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"FE32")

      port map(A => \sercon_8_0_2[3]\, B => un5_penable, C => 
        N_161, D => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \sercon_9[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => \fsmsta[18]_net_1\, B => N_2177, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \serdat_RNIE9801[7]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(7), B => \serdat[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_RNO\ : CFG3
      generic map(INIT => x"8C")

      port map(A => N_2177, B => N_191, C => \un151_framesync\, Y
         => N_193);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un1_ens1\ : CFG2
      generic map(INIT => x"4")

      port map(A => \adrcomp\, B => \fsmmod[6]_net_1\, Y => 
        un1_ens1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2171, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6s2\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sm0);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3_0[19]\ : CFG4
      generic map(INIT => x"001F")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \SDAInt\, D => N_2177, Y => \fsmsta_8_i_a3_0[19]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \sercon[6]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \un1_PCLK_count1_1.CO0\ : CFG3
      generic map(INIT => x"40")

      port map(A => \PCLK_count1_ov_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1[0]_net_1\, Y => 
        CO0_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"D555")

      port map(A => N_2176, B => N_2187, C => N_95, D => 
        \adrcomp_2_sqmuxa_i_a3_4\, Y => adrcomp_2_sqmuxa_i_0_5);
    
    \un2_framesync_1_1.CO1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CO0, B => \framesync[1]_net_1\, Y => CO1_2);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"02")

      port map(A => N_1656, B => fsmsta_8_23_351_i_0_1, C => 
        N_2181, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \fsmsync_ns_0_a3_2_2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[4]_net_1\, Y
         => N_1002_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG4
      generic map(INIT => x"0045")

      port map(A => \adrcomp\, B => \framesync[0]_net_1\, C => 
        \framesync[3]_net_1\, D => \fsmsta_cnst[0]\, Y => 
        fsmsta_8_9_509_0_1);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0045")

      port map(A => bsd7_9_iv_1, B => \serdat[7]_net_1\, C => 
        bsd7_tmp_6_sn_N_10_mux, D => bsd7_i_m, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \indelay[1]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_6[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[15]_net_1\, 
        C => un135_ens1_2, Y => \sersta_32_6[2]\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \sersta_RNIAV3U1[3]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        seradr0apb(6), Y => N_1220);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.ANC2\ : CFG3
      generic map(INIT => x"07")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[2]_net_1\, Y
         => ANC2);
    
    \serSTA_WRITE_PROC.sersta_32_5[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[24]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[0]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_5[2]\);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(3), B => seradr0apb(2), C => 
        \serdat[2]_net_1\, D => \serdat[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    adrcomp_2_sqmuxa_i_a3_1 : CFG2
      generic map(INIT => x"8")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, Y => \adrcomp_2_sqmuxa_i_a3_1\);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_11_454_i_a6_2_0_0_o2\ : CFG3
      generic map(INIT => x"DF")

      port map(A => \adrcomp\, B => \fsmsta[23]_net_1\, C => 
        \adrcompen\, Y => N_2182);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_2, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"515F")

      port map(A => \fsmsta[11]_net_1\, B => N_2186, C => N_2177, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[0]_net_1\, C
         => \fsmsta[5]_net_1\, D => \fsmsta[4]_net_1\, Y => 
        \sersta_32_i_a2_9[3]\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[1]_net_1\, C
         => \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => N_2177, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, Y
         => N_629);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_6_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \fsmmod_ns_0_a4_0_1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \starto_en\, B => N_64, C => N_1040, D => 
        un115_fsmdet, Y => N_1059_1);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    un1_fsmsta_1_i_0_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[12]_net_1\, 
        C => \fsmsta[16]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => N_1470, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => un135_ens1_7, B => \fsmsta[14]_net_1\, Y => 
        N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \serCON_WRITE_PROC.un3_penable_0_0\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), B => 
        CoreAPB3_0_APBmslave0_PWRITE, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), D => 
        CoreAPB3_0_APBmslave0_PENABLE, Y => un3_penable_0);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    SDAO_int_RNI3J14 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_6_SDAO[0]\, Y => 
        COREI2C_0_6_SDAO_i(0));
    
    \sersta_RNI6R3U1[2]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        \sercon[5]_net_1\, Y => N_1219);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[26]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_18_s5_1_0, Y => 
        \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG3
      generic map(INIT => x"21")

      port map(A => \framesync[3]_net_1\, B => N_92, C => 
        \framesync[0]_net_1\, Y => un74_ens1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[21]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"8C00")

      port map(A => \framesync[3]_net_1\, B => N_1717, C => 
        N_1652, D => fsmsta_8_3_601_0_1, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_ns_0_a4[5]\ : CFG3
      generic map(INIT => x"04")

      port map(A => un115_fsmdet, B => \fsmmod[1]_net_1\, C => 
        un10_sclscl, Y => N_1058);
    
    PCLK_count1_1_sqmuxa_0 : CFG4
      generic map(INIT => x"002F")

      port map(A => \PCLK_count1[2]_net_1\, B => CO1_0, C => 
        \PCLK_count1_0_sqmuxa_4_1\, D => \PCLK_count1_0_sqmuxa_3\, 
        Y => \PCLK_count1_1_sqmuxa_0\);
    
    \fsmmod_ns_0_a4[0]\ : CFG4
      generic map(INIT => x"AAA2")

      port map(A => \fsmmod[6]_net_1\, B => \starto_en\, C => 
        N_1040, D => N_64, Y => N_1048);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \sersta_32_i_a2_8[4]\, B => 
        \sersta_32_i_a2_6[4]\, C => \sersta_32_i_a2_7[4]\, D => 
        \sersta_32_i_a2_5[4]\, Y => N_100_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"C5")

      port map(A => N_2196, B => \COREI2C_0_6_SDAO[0]\, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \ack\, B => N_2177, C => N_133, D => 
        fsmsta_8_28_307_a3_0_1, Y => N_1486);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"27")

      port map(A => un33_fsmsta, B => \nedetect\, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG3
      generic map(INIT => x"20")

      port map(A => \PCLK_count1_1_sqmuxa_4\, B => 
        \PCLK_count1_ov_1_sqmuxa\, C => PCLK_count2_ov_6_1, Y => 
        \PCLK_count1_1_sqmuxa\);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serdat_RNIJ7T11[4]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[4]_net_1\, B => \sercon[4]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[4]\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[6]_net_1\, C
         => \fsmmod[1]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"02")

      port map(A => N_2196, B => \COREI2C_0_6_SDAO[0]\, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \un1_counter_rst_3\, D => 
        CO0_0, Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => \fsmsta[16]_net_1\, B => N_2177, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_1, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \sersta_RNIE34U1[4]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        \sercon[7]_net_1\, Y => N_1221);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"00D0")

      port map(A => N_2186, B => N_2177, C => N_82, D => 
        un136_framesync, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"88A8")

      port map(A => \SCLInt\, B => \fsmdet[3]_net_1\, C => 
        \fsmdet[2]_net_1\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \sersta_32_4[1]\, B => m7_3, C => 
        \sersta_32_5[1]\, D => m7_4, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[27]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_24_s4_1_0, Y => 
        \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[3]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmsta[21]_net_1\, B => \fsmsta[22]_net_1\, 
        C => \COREI2C_0_6_INT[0]\, Y => \sersta_32_i_a2_6[3]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[3]\ : CFG4
      generic map(INIT => x"7F80")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, C => CO0, D => \framesync[3]_net_1\, 
        Y => \framesync_7_enl_bm_2[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG4
      generic map(INIT => x"3600")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => N_92, D => N_2179, Y => 
        N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG3
      generic map(INIT => x"54")

      port map(A => N_2181, B => fsmsta_8_5_555_a3_0_2, C => 
        fsmsta_8_5_555_a3_2, Y => N_1665);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    PCLKint_ff_RNIRBPH : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_6_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"7075")

      port map(A => \ack\, B => un13_adrcompen, C => 
        \adrcomp_2_sqmuxa_i_a2_1_5\, D => N_133, Y => N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_6_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => N_1470);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    PCLK_count1_0_sqmuxa_4_1 : CFG3
      generic map(INIT => x"01")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \PCLK_count1_0_sqmuxa_4_1\);
    
    PCLK_count1_1_sqmuxa_1_0 : CFG4
      generic map(INIT => x"CCFA")

      port map(A => \sercon[1]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \sercon[7]_net_1\, D => 
        \PCLK_count1_1_sqmuxa_1_0_1\, Y => 
        \PCLK_count1_1_sqmuxa_1_0\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \fsmsta_RNO[19]\ : CFG4
      generic map(INIT => x"000B")

      port map(A => N_191, B => \fsmsta_8_i_a3_0[19]\, C => 
        N_2199, D => un136_framesync, Y => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_92, B => \framesync[0]_net_1\, Y => N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \COREI2C_0_6_INT[0]\, B => \sercon[5]_net_1\, 
        C => N_1041, D => \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => 
        N_1054);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_0\ : CFG4
      generic map(INIT => x"F3FA")

      port map(A => N_2182, B => \fsmsta[9]_net_1\, C => N_2181, 
        D => N_2177, Y => fsmsta_8_4_577_i_0);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_0_2\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[4]_net_1\, Y => fsmsta_8_9_509_a4_0);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[12]_net_1\, 
        C => \fsmsta[22]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        un25_fsmsta_1);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFBA")

      port map(A => un16_fsmmod, B => N_2177, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_6_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \fsmmod_ns_i_o3_1_1[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, Y => N_92);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO0, B => framesync_7_e2, C => 
        \framesync[1]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[1]\);
    
    \sersta_RNIUI3U1[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => un16_fsmmod, B => \sercon_8_2[4]\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), D => un5_penable, Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => N_76, D => \fsmsync[4]_net_1\, Y => N_55_i_0);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG4
      generic map(INIT => x"AEAA")

      port map(A => N_2181, B => un91_ens1, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"8090")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1_ov_1_sqmuxa\, C => PCLK_count2_ov_6_1, D => 
        \PCLK_count1_1_sqmuxa_4\, Y => \PCLK_count1_10[0]\);
    
    \serSTA_WRITE_PROC.sersta_32_4[0]\ : CFG4
      generic map(INIT => x"FEFF")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, C
         => \fsmsta[9]_net_1\, D => \COREI2C_0_6_INT[0]\, Y => 
        \sersta_32_4[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, Y => 
        un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO\ : CFG4
      generic map(INIT => x"C010")

      port map(A => \nedetect\, B => \COREI2C_0_6_INT[0]\, C => 
        bsd7_i_m_0, D => un105_ens1, Y => bsd7_i_m);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, C
         => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[0]\ : CFG4
      generic map(INIT => x"07FF")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_e2_1, Y => 
        \framesync_7_enl_am[0]\);
    
    \fsmmod_ns_0_a4[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \nedetect\, B => un115_fsmdet, C => 
        \fsmmod[5]_net_1\, Y => N_1050);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    \un2_framesync_1_1.CO0\ : CFG4
      generic map(INIT => x"8808")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync[3]_net_1\, D => N_92, Y => CO0);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"22EF")

      port map(A => \COREI2C_0_6_SDAO[0]\, B => N_2177, C => 
        \fsmsta[22]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"3031")

      port map(A => N_1041, B => N_1043, C => \fsmmod[2]_net_1\, 
        D => N_997, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un3_penable_0, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), C => 
        N_8_0, D => un5_penable_1, Y => un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    PCLK_count1_0_sqmuxa_2 : CFG4
      generic map(INIT => x"0545")

      port map(A => \sercon[7]_net_1\, B => CO1, C => 
        \PCLK_count1[3]_net_1\, D => \PCLK_count1[2]_net_1\, Y
         => \PCLK_count1_0_sqmuxa_2\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG3
      generic map(INIT => x"20")

      port map(A => un137_framesync, B => \ack\, C => 
        un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => \sercon[5]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"4440")

      port map(A => un16_fsmmod, B => PCLK_count2_ov_6_0_a2_1_3, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    un1_counter_rst_3 : CFG3
      generic map(INIT => x"5D")

      port map(A => PCLK_count2_ov_6_1, B => 
        \PCLK_count1_1_sqmuxa_4\, C => \PCLK_count1_ov_1_sqmuxa\, 
        Y => \un1_counter_rst_3\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta[5]_net_1\, C
         => \fsmsta[4]_net_1\, D => \fsmsta[13]_net_1\, Y => 
        \sersta_32_i_a2_8[4]\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_6_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, C => \framesync[3]_net_1\, D => 
        \framesync[0]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"ACAA")

      port map(A => \fsmsta[13]_net_1\, B => 
        \COREI2C_0_6_SDAO[0]\, C => N_2177, D => N_2196, Y => 
        N_82);
    
    \fsmsta_RNO[12]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => N_2181, B => N_1656, C => N_2186, D => N_124, 
        Y => N_1774_i_0);
    
    PCLK_count1_ov_1_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \sercon[7]_net_1\, B => bclke, C => 
        \sercon[1]_net_1\, D => \sercon[0]_net_1\, Y => 
        \PCLK_count1_ov_1_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_6_SDAO[0]\, Y => 
        N_172);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_m1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un92_fsmsta, Y => bsd7_tmp_6_m1);
    
    adrcomp : SLE
      port map(D => N_2176, CLK => FAB_CCC_GL0, EN => 
        adrcomp_2_sqmuxa_i_0_5, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[11]_net_1\, C
         => \fsmsta[7]_net_1\, D => \fsmsta[23]_net_1\, Y => m7_4);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \fsmdet[3]_net_1\, B => N_629, C => 
        \fsmdet[1]_net_1\, Y => N_1717);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_5\ : CFG2
      generic map(INIT => x"E")

      port map(A => un135_ens1_2, B => un135_ens1_7, Y => 
        un135_ens1_5);
    
    un1_fsmsta_i_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[18]_net_1\, 
        Y => un135_ens1_7);
    
    \serCON_WRITE_PROC.un91_ens1_0_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \pedetect\, Y => un91_ens1);
    
    \fsmmod_RNI0I621[5]\ : CFG4
      generic map(INIT => x"FEF0")

      port map(A => \fsmmod[0]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmsta_cnst[0]\, D => \fsmdet[3]_net_1\, Y => 
        N_1622_2);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \fsmsta[9]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \PCLKint\, B => \PCLKint_ff\, C => N_1586_1, 
        D => \fsmmod[2]_net_1\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1041, B => N_997, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[26]\);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => N_1665, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \fsmsync[5]_net_1\, B => N_64, C => 
        \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0_o4[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => un115_fsmdet, B => N_1064, Y => N_1043);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_RNIU1491\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \nedetect\, B => \COREI2C_0_6_INT[0]\, C => 
        un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sn_N_10_mux);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1050, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_6_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => un135_ens1_2, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_2181, B => N_1656, C => 
        fsmsta_8_2_647_i_0_0, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_3\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[8]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[16]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[22]\, B => un136_framesync, C
         => \fsmsta[22]_net_1\, D => N_2177, Y => \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_5, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \framesync_7_enl_bm[0]\, B => 
        \framesync_7_enl_am[0]\, C => framesync_7_e2, Y => 
        \framesync_7[0]\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG3
      generic map(INIT => x"06")

      port map(A => \PCLK_count1[1]_net_1\, B => CO0_0, C => 
        \un1_counter_rst_3\, Y => \PCLK_count1_10[1]\);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_64, D => N_1002_3, Y => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \bsd7_tmp\, B => \SCLInt\, C => 
        \COREI2C_0_6_INT[0]\, D => un57_fsmsta, Y => 
        bsd7_tmp_i_m_2);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"F0F8")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat_2_sqmuxa_1_0\, Y => 
        un1_serdat_2_sqmuxa_5);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serdat_RNINBT11[6]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[6]_net_1\, B => \sercon[6]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1002, B => \COREI2C_0_6_INT[0]\, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_6_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_6_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"0C08")

      port map(A => un92_fsmsta, B => \pedetect\, C => un105_ens1, 
        D => \un1_serdat40\, Y => \un1_serdat_2_sqmuxa_1\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_7\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, D => un135_ens1_5, Y => 
        un135_ens1_7_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_26_328_a3_0_1_i\ : CFG2
      generic map(INIT => x"7")

      port map(A => \fsmsta[23]_net_1\, B => \adrcomp\, Y => N_26);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_6\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[23]_net_1\, C
         => fsmsta_8_20_379_i_0_a3_3_0, D => 
        fsmsta_8_20_379_i_0_a3_4, Y => fsmsta_8_20_379_i_0_a3_6);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[3]_net_1\, B => \fsmsta[13]_net_1\, C
         => \fsmsta[23]_net_1\, Y => \adrcomp_2_sqmuxa_i_o2_1_2\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_3_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF20")

      port map(A => fsmsta_8_3_601_a4_0, B => \fsmdet[1]_net_1\, 
        C => N_1656, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_172, B => N_2193, C => N_2182, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_1002_3, B => 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[2]_net_1\, Y => N_1002);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[27]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[3]_net_1\, B => \serdat[2]_net_1\, C
         => \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[26]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \ack\, B => \adrcompen\, C => N_2177, D => 
        N_26, Y => fsmsta_8_5_555_a3_0_2);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_6_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3340")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => un1_fsmmod, D => N_1586_1, Y => N_1624);
    
    adrcomp_2_sqmuxa_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[23]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => N_95);
    
    PCLK_count1_1_sqmuxa_1_0_1 : CFG4
      generic map(INIT => x"1808")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => CO1, D => bclke, Y => 
        \PCLK_count1_1_sqmuxa_1_0_1\);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_6_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        \COREI2C_0_6_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a4_0_3\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmsta[10]_net_1\, Y => fsmsta_8_3_601_a4_0);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_1046, B => N_1054, C => 
        \fsmmod_ns_i_0[2]_net_1\, D => un115_fsmdet, Y => 
        N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNI7FEF : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        un136_framesync, C => \pedetect\, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \serCON_WRITE_PROC.sercon_8_0_1[3]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \sercon[6]_net_1\, B => N_2179, C => 
        un91_ens1, D => N_163, Y => \sercon_8_0_1[3]\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[6]_net_1\, B => \fsmsync[3]_net_1\, 
        C => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_1, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \sersta_RNI2N3U1[1]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[4]\, C => \sersta[1]_net_1\, D => 
        seradr0apb(4), Y => N_1218);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    \fsmsync_ns_i_1[6]\ : CFG4
      generic map(INIT => x"F7F4")

      port map(A => \SDAInt\, B => \fsmsync[1]_net_1\, C => 
        N_1002, D => N_997, Y => \fsmsync_ns_i_1[6]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => N_1449, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_6_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[16]_net_1\, 
        C => \fsmsta[19]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5\ : CFG4
      generic map(INIT => x"0400")

      port map(A => un1_fsmmod, B => N_1466, C => 
        \fsmmod[2]_net_1\, D => N_629, Y => N_1467);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => N_2177, B => fsmsta_8_20_379_i_0_a3_6, C => 
        N_2181, D => N_91, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"3100")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_e2_1, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[6]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \CLK_COUNTER1_PROC.un12_pclk_count1_1.ANC1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \PCLK_count1[0]_net_1\, Y => CO1);
    
    \FSMSTA_SYNC_PROC.un137_framesync\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un91_ens1, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => un137_framesync);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \fsmsync_ns_i_a3_1_0_a2_1[2]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, Y
         => \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"8C00")

      port map(A => \framesync[3]_net_1\, B => N_1717, C => 
        N_1652, D => fsmsta_8_9_509_0_1, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_126, B => N_80, C => un136_framesync, Y => 
        N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"FBF8")

      port map(A => \PWDATA_i_m_1[7]\, B => un105_ens1, C => 
        \fsmdet[3]_net_1\, D => bsd7_tmp_i_m_2, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \PCLKint\, B => \un151_framesync\, C => 
        \PCLKint_ff\, Y => \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \fsmsync_ns_i_o3_0[6]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => un70_fsmsta, B => \fsmsync[5]_net_1\, C => 
        N_64, Y => N_995);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[9]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF20")

      port map(A => fsmsta_8_9_509_a4_0, B => \fsmdet[1]_net_1\, 
        C => N_1656, D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"5444")

      port map(A => un115_fsmdet, B => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, C => \fsmmod[3]_net_1\, D
         => N_1034, Y => \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FDFF")

      port map(A => m7_3, B => \sersta_32_3[0]\, C => 
        \sersta_32_4[0]\, D => m7_4, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        C => un135_ens1_7_0, D => un135_ens1_3, Y => un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_5, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[0]_net_1\, C
         => un1_ens1, Y => \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    un1_serdat_2_sqmuxa_1_0 : CFG4
      generic map(INIT => x"00EF")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => un57_fsmsta, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1_0\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => \bsd7_tmp\, B => bsd7_tmp_6_m1, C => 
        bsd7_tmp_6_sm0, D => bsd7_tmp_6_sn_N_10_mux, Y => 
        bsd7_tmp_6);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un3_penable_0, B => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), C => 
        N_8_0, D => un105_ens1_1, Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"3100")

      port map(A => un74_ens1, B => N_1622_2, C => 
        \COREI2C_0_6_INT[0]\, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0_RNIVEM21\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => un57_fsmsta_1_0, Y => N_191);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \fsmsync_RNO[1]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => N_995, B => \fsmsync_ns_i_1[6]_net_1\, C => 
        \fsmsync[1]_net_1\, D => \fsmsync[2]_net_1\, Y => 
        N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1058, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => \fsmsta[28]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \serCON_WRITE_PROC.sercon_8_0_2[3]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \sercon[6]_net_1\, B => \COREI2C_0_6_INT[0]\, 
        C => \sercon_8_0_1[3]\, D => N_134, Y => 
        \sercon_8_0_2[3]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_6_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[3]\ : CFG4
      generic map(INIT => x"07FF")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_e2_1, Y => 
        \framesync_7_enl_am_2[3]\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[4]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmsta[6]_net_1\, B => \fsmsta[14]_net_1\, C
         => \COREI2C_0_6_INT[0]\, Y => \sersta_32_i_a2_5[4]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[5]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG4
      generic map(INIT => x"0307")

      port map(A => \fsmmod[0]_net_1\, B => \nedetect\, C => 
        \fsmmod[4]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \fsmmod_ns_i_0[2]_net_1\);
    
    \FSMMOD_COMB_PROC.un10_sclscl\ : CFG2
      generic map(INIT => x"8")

      port map(A => \pedetect\, B => \SCLSCL\, Y => un10_sclscl);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_1586_1, B => N_2177, C => \fsmsta[8]_net_1\, 
        D => N_172, Y => fsmsta_8_5_555_a3_2);
    
    \fsmmod_ns_i_o3_0_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_6_INT[0]\, B => \sercon[4]_net_1\, 
        Y => N_997);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    SCLO_int_RNID421 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_6_SCLO[0]\, Y => 
        COREI2C_0_6_SCLO_i(0));
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1_3, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG3
      generic map(INIT => x"02")

      port map(A => un137_framesync, B => \ack\, C => 
        un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_5);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmdet[3]_net_1\, B => un139_ens1_0, C => 
        \fsmdet[1]_net_1\, Y => framesync_7_e2_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_5 is

    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          COREI2C_0_6_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 2);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 12);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          un3_penable                                : in    std_logic;
          bclke                                      : in    std_logic;
          N_1218                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          BIBUF_COREI2C_0_6_SCL_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_6_SDA_IO_Y                 : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_8_0                                      : in    std_logic;
          un105_ens1_1                               : in    std_logic;
          un5_penable_1                              : in    std_logic
        );

end COREI2C_5;

architecture DEF_ARCH of COREI2C_5 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_5
    port( COREI2C_0_6_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 2) := (others => 'U');
          seradr0apb                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          bclke                                      : in    std_logic := 'U';
          N_1218                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          BIBUF_COREI2C_0_6_SCL_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_6_SDA_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_8_0                                      : in    std_logic := 'U';
          un105_ens1_1                               : in    std_logic := 'U';
          un5_penable_1                              : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_5
	Use entity work.COREI2CREAL_6_5(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_5
      port map(COREI2C_0_6_SDAO_i(0) => COREI2C_0_6_SDAO_i(0), 
        COREI2C_0_6_SCLO_i(0) => COREI2C_0_6_SCLO_i(0), 
        COREI2C_0_6_INT(0) => COREI2C_0_6_INT(0), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, bclke => bclke, N_1218 => 
        N_1218, N_1221 => N_1221, N_1219 => N_1219, N_1217 => 
        N_1217, N_1220 => N_1220, BIBUF_COREI2C_0_6_SCL_IO_Y => 
        BIBUF_COREI2C_0_6_SCL_IO_Y, BIBUF_COREI2C_0_6_SDA_IO_Y
         => BIBUF_COREI2C_0_6_SDA_IO_Y, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, N_8_0 => N_8_0, 
        un105_ens1_1 => un105_ens1_1, un5_penable_1 => 
        un5_penable_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_3 is

    port( COREI2C_0_4_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_INT                            : out   std_logic_vector(0 to 0);
          seradr0apb                                 : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 1);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 13);
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          BIBUF_COREI2C_0_4_SDA_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_4_SCL_IO_Y                 : in    std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic;
          un3_penable_1                              : in    std_logic;
          un105_ens1_3                               : in    std_logic;
          un5_penable_2                              : out   std_logic;
          bclke                                      : in    std_logic;
          N_8_0                                      : in    std_logic;
          N_43                                       : in    std_logic;
          un105_ens1_0                               : in    std_logic
        );

end COREI2CREAL_6_3;

architecture DEF_ARCH of COREI2CREAL_6_3 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_4_SDAO[0]\, \COREI2C_0_4_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_4_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        un1_serdat_2_sqmuxa_3, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, N_1665, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, N_1470, \ack\, ack_7, 
        SDAO_int_7_0_275, SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, 
        bsd7_tmp_6, \bsd7\, bsd7_9_iv_i_0, \adrcomp\, N_2176, 
        adrcomp_2_sqmuxa_i_0_3, \PCLKint\, PCLKint_3, 
        un1_pclkint4_i_0, \ack_bit\, \ack_bit_1_sqmuxa\, 
        \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_3, un1_rtn_3_3, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, PCLK_count2_ov_6_1, 
        \un1_PCLK_count1_0_sqmuxa\, CO1, N_126, N_2181, 
        un133_framesync, N_80, un57_fsmsta, \un1_serdat40\, 
        \un1_serdat_2_sqmuxa_1_0\, un91_ens1, 
        \adrcomp_2_sqmuxa_i_o2_1_3\, \un1_fsmsta_1_i_0_o2_0\, 
        un25_fsmsta_1, un25_fsmsta, un16_fsmmod, \sersta_32_5[2]\, 
        N_1586_1, un105_ens1, N_2177, N_2173_i_1, N_133, 
        un1_fsmmod, N_36_i_1, un136_framesync, N_2196, N_2186, 
        \un1_PCLK_count1_0_sqmuxa_1\, 
        \un1_PCLK_count1_0_sqmuxa_0\, 
        \un1_PCLK_count1_0_sqmuxa_1_0\, CO2, ANC2, 
        \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, 
        \fsmsta_cnst[0]\, fsmsta_8_9_509_0_1, N_1717, 
        fsmsta_8_9_509_0, N_1652, fsmsta_8_3_601_0_1, 
        fsmsta_8_3_601_0, \un1_pclk_count1_ov_1_1\, 
        \un1_pclk_count1_ov_1\, un135_ens1_1, un135_ens1_7, 
        un135_ens1_2, un135_ens1, \adrcomp_2_sqmuxa_i_o2_1_1\, 
        un135_ens1_3, \PRDATA_3_1[4]\, \PRDATA_3_1_1[5]\, 
        \PRDATA_3_1[3]\, \PRDATA_3_1_1[6]\, \PRDATA_3_1_1[7]\, 
        \fsmsta_8_ns_1[18]\, un13_adrcompen, \fsmsta_8_ns_1[28]\, 
        \fsmsta_8_ns_1[29]\, \fsmsta_8_ns_1[16]\, framesync_7_e2, 
        \framesync_7_enl_bm_0[3]\, \framesync_7_enl_am_0[3]\, 
        \framesync_7_enl_bm_0[0]\, \framesync_7_enl_am_0[0]\, 
        N_2179, N_161_2, PCLK_count2_ov_6_0_a2_1_0, 
        un111_fsmdet_0, \sersta_32_i_a2_5[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, un139_ens1_0, N_67, 
        mst, un26_adrcompen_6, N_145_2, N_23, N_127, N_64, 
        N_1002_3, \un151_framesync\, N_1196, N_1197, N_1198, 
        SDAO_int_7_0_275_1, \adrcomp_2_sqmuxa_i_a3_3\, 
        SDAO_int_7_0_275_a5_0, un141_ens1_2, 
        \SDAO_int_1_sqmuxa_3\, \adrcomp_2_sqmuxa_i_a2_1_2\, 
        \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_5_555_a3_0_1, 
        fsmsta_8_10_476_i_a6_1, fsmsta_8_5_555_a3_0, 
        \fsmmod_ns_i_a4_1_0[2]_net_1\, \sersta_32_5[1]\, 
        \sersta_32_4[1]\, \sersta_32_4[0]\, \sersta_32_3[0]\, 
        fsmsta_8_20_379_i_0_a3_5, fsmsta_8_20_379_i_0_a3_4, 
        \sersta_32_i_a2_7[4]\, \sersta_32_i_a2_6[4]\, 
        \sersta_32_4[2]\, fsmsta_nxt_1_sqmuxa_24_s4_1_0, 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0, \sersta_32_i_a2_8[3]\, 
        \sersta_32_i_a2_7[3]\, un13_adrcompen_4, m7_5, m7_4, 
        \PCLK_count1_ov_1_sqmuxa_1\, un12_pclk_count1, N_1064, 
        un33_fsmsta, framesync_7_sm0, 
        PCLK_count2_ov_6_0_a2_1_4_tz, N_1034, N_68, CO1_0, N_76, 
        CO2_0, \un1_pclk_count1_ov\, N_1049, N_163_2, N_189, N_95, 
        un70_fsmsta, N_2182, N_1040, \adrcomp_2_sqmuxa_i_a3_4\, 
        \fsmmod_ns_i_0[2]_net_1\, fsmsta_8_10_476_i_0, 
        \SDAO_int_1_sqmuxa_4\, \fsmsync_ns_i_0[6]_net_1\, 
        \adrcomp_2_sqmuxa_i_a2_1_4\, PCLK_count2_ov_6_0_a2_1_3, 
        \fsmsta_8_i_a3_0[19]\, \sersta_32_i_a2_9[4]\, 
        \sercon_8_2[4]\, \sersta_32_7[2]\, \sersta_32_i_a2_10[3]\, 
        N_1002, N_104, \PCLK_count1_0_sqmuxa_4\, N_2192, 
        un19_framesync, un25_framesync, \fsmsta_8_0_a2_1[7]\, 
        N_130, N_63, N_84, \un1_pclk_count191\, N_1622_2, N_1732, 
        N_2171, N_2193, N_191, \un1_fsmsta_6\, un74_ens1, N_1041, 
        N_1656, N_120, N_124, fsmsta_8_28_307_a3_0_1, 
        \SDAO_int_1_sqmuxa_7\, \adrcomp_2_sqmuxa_i_a2_1_5\, 
        N_1007, N_162, N_165, \fsmsta_nxt_9_m[27]\, 
        \fsmsta_nxt_9_m[26]\, \fsmsta_nxt_9_m[21]\, 
        \fsmsta_nxt_9_m[22]\, N_1054, un115_fsmdet, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, \un5_penable_2\, N_1046, 
        \PCLK_count1_0_sqmuxa_3\, N_1624, N_1657_2, N_70, CO0, 
        N_1060, N_1048, \fsmsta_8_i_0[25]\, fsmsta_8_4_577_i_0, 
        N_82, bsd7_i_m_0, bsd7_tmp_i_m_2, 
        fsmsta_8_20_379_i_0_o2_0, \sercon_8_0_1[3]\, 
        \sercon_8_0_0[3]\, \fsmsync_ns_0_0_1[0]_net_1\, 
        fsmsta_8_23_351_i_0_1, \un1_ens1_pre_1_sqmuxa_0_a2_1\, 
        N_1465, N_1680, N_145, N_166, N_1058, N_1050, 
        \fsmsync_ns_i_0_1_tz[3]_net_1\, N_86, un92_fsmsta, 
        un1_fsmsta_10_i_0, CO1_1, N_1059_1, N_2199, 
        \PWDATA_i_m_1[7]\, fsmsta_8_2_647_i_0_0, N_1486, 
        un134_fsmsta, \serdat_0_sqmuxa\, N_2187, N_1466, 
        bsd7_tmp_6_sn_N_10_mux, \sercon_8[3]\, bsd7_tmp_6_m1, 
        bsd7_tmp_6_sm0, bsd7_9_iv_1, \un1_counter_rst_3\, 
        bsd7_i_m, \un1_serdat_2_sqmuxa_1\ : std_logic;

begin 

    COREI2C_0_4_INT(0) <= \COREI2C_0_4_INT[0]\;
    un5_penable_2 <= \un5_penable_2\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    adrcomp_2_sqmuxa_i_0_0 : CFG4
      generic map(INIT => x"0015")

      port map(A => un16_fsmmod, B => N_2192, C => 
        \COREI2C_0_4_INT[0]\, D => N_1586_1, Y => N_2176);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmmod_RNIKNAQ[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_189, B => \fsmsta_cnst[0]\, Y => N_1622_2);
    
    \fsmsync_ns_i_a3_0[6]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[1]_net_1\, 
        C => N_68, D => un70_fsmsta, Y => N_1007);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[0]_net_1\, B => seradr0apb(1), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_145_2, 
        Y => N_2171);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_191, B => \un1_fsmsta_6\, C => 
        \fsmsta[23]_net_1\, D => un1_fsmmod, Y => N_166);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => framesync_7_e2, B => 
        \framesync_7_enl_bm_0[3]\, C => \framesync_7_enl_am_0[3]\, 
        Y => \framesync_7[3]\);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \adrcomp_2_sqmuxa_i_o2_1_1\, 
        Y => un19_framesync);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[2]_net_1\, B => seradr0apb(3), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_6, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_3, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \bsd7\, Y => bsd7_i_m_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[0]\ : CFG3
      generic map(INIT => x"36")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        un70_fsmsta, Y => \framesync_7_enl_bm_0[0]\);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_1656, B => \fsmdet[1]_net_1\, Y => N_1657_2);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => \un1_fsmsta_1_i_0_o2_0\, D => un25_fsmsta_1, Y => 
        un25_fsmsta);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sersta_32_5[2]\, B => \sersta_32_7[2]\, C
         => un135_ens1_2, D => \un1_fsmsta_1_i_0_o2_0\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1041, B => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, 
        C => N_1040, Y => \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    \fsmmod_ns_0[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_1064, B => N_1049, C => un115_fsmdet, D => 
        N_1048, Y => \fsmmod_ns[0]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_1\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => N_2181, C => 
        \adrcompen\, D => \adrcomp\, Y => fsmsta_8_28_307_a3_0_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => un1_fsmmod, B => SDAO_int_7_0_275_a5_0, C => 
        N_1466, D => SDAO_int_7_0_275_1, Y => SDAO_int_7_0_275);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[2]_net_1\);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \sercon[7]_net_1\, D => 
        \un1_pclk_count1_ov_1_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => un139_ens1_0, Y => 
        framesync_7_sm0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"003A")

      port map(A => \ack\, B => N_172, C => N_2177, D => 
        fsmsta_8_4_577_i_0, Y => N_2172_i_0);
    
    \fsmmod_ns_0_a4_0[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[1]_net_1\, B => \SCLSCL\, C => 
        \pedetect\, Y => N_1049);
    
    un1_PCLK_count1_0_sqmuxa_0 : CFG4
      generic map(INIT => x"FF10")

      port map(A => \sercon[1]_net_1\, B => \sercon[7]_net_1\, C
         => un12_pclk_count1, D => \PCLK_count1_0_sqmuxa_4\, Y
         => \un1_PCLK_count1_0_sqmuxa_0\);
    
    \fsmsta_RNO[25]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => N_172, B => N_2177, C => \fsmsta_8_i_0[25]\, 
        D => un136_framesync, Y => N_2175_i_0);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_6\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), Y => 
        un26_adrcompen_6);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync[2]_net_1\, D => \framesync[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \fsmsta[17]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1652, D => un1_fsmmod, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_3_601_0_1);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_4_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1586_1, B => \fsmsta[8]_net_1\, Y => 
        fsmsta_8_5_555_a3_0);
    
    \un1_PCLK_count1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \un1_PCLK_count1_0_sqmuxa\, C => \PCLK_count1[1]_net_1\, 
        Y => CO1);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"F780")

      port map(A => \un5_penable_2\, B => N_43, C => 
        CoreAPB3_0_APBmslave0_PWDATA(3), D => \sercon_8[3]\, Y
         => \sercon_9[3]\);
    
    PCLK_count1_0_sqmuxa_4 : CFG4
      generic map(INIT => x"0004")

      port map(A => \sercon[7]_net_1\, B => CO2_0, C => 
        \sercon[1]_net_1\, D => \sercon[0]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[18]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.CO2\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2_0);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_3);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6s2\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sm0);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[7]_net_1\);
    
    PCLK_count1_ov_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \PCLK_count1_ov_1_sqmuxa_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3_0[19]\ : CFG4
      generic map(INIT => x"001F")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \SDAInt\, D => N_2177, Y => \fsmsta_8_i_a3_0[19]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => mst, D => \sercon[6]_net_1\, Y => \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"D555")

      port map(A => N_2176, B => N_2187, C => 
        \adrcomp_2_sqmuxa_i_a3_4\, D => N_95, Y => 
        adrcomp_2_sqmuxa_i_0_3);
    
    \un2_framesync_1_1.CO1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CO0, B => \framesync[1]_net_1\, Y => CO1_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[2]_net_1\, C
         => \fsmmod[0]_net_1\, Y => SDAO_int_7_0_275_a5_0);
    
    un151_framesync : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        Y => \un151_framesync\);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"10")

      port map(A => fsmsta_8_23_351_i_0_1, B => N_2181, C => 
        N_1656, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \fsmsync_ns_0_a3_2_2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[4]_net_1\, Y
         => N_1002_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_9_509_0_1);
    
    \serCON_WRITE_PROC.sercon_8_0[3]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => N_161_2, B => \sercon_8_0_1[3]\, C => N_163_2, 
        D => \sercon_8_0_0[3]\, Y => \sercon_8[3]\);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0045")

      port map(A => bsd7_9_iv_1, B => \serdat[7]_net_1\, C => 
        bsd7_tmp_6_sn_N_10_mux, D => bsd7_i_m, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \indelay[1]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.ANC2\ : CFG3
      generic map(INIT => x"15")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => ANC2);
    
    \serSTA_WRITE_PROC.sersta_32_5[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[24]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_5[2]\);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(4), B => seradr0apb(2), C => 
        \serdat[3]_net_1\, D => \serdat[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a3_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta_cnst[0]\, B => \fsmdet[3]_net_1\, Y
         => N_1732);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_11_454_i_a6_2_0_0_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, Y => 
        N_2182);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO1_1, B => framesync_7_e2, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"4577")

      port map(A => \fsmsta[11]_net_1\, B => N_2177, C => N_2186, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[2]_net_1\, C
         => \fsmsta[12]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \fsmmod_RNIV7TC[5]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmdet[3]_net_1\, Y => N_189);
    
    \serdat_RNILPIV[7]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[7]_net_1\, B => \sercon[7]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => N_2177, Y => N_2193);
    
    \serdat_RNI2RB11[3]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(3), B => \serdat[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1[3]\);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_4_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \fsmmod_ns_0_a4_0_1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \starto_en\, B => N_64, C => N_1040, D => 
        un115_fsmdet, Y => N_1059_1);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    un1_fsmsta_1_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => 
        \fsmsta[12]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => N_1470, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => un135_ens1_7, B => \fsmsta[14]_net_1\, Y => 
        N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_1[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1586_1, B => \sercon[6]_net_1\, Y => 
        N_163_2);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_0\ : CFG4
      generic map(INIT => x"C055")

      port map(A => \fsmsta[3]_net_1\, B => \framesync[0]_net_1\, 
        C => \framesync[3]_net_1\, D => N_1586_1, Y => 
        fsmsta_8_10_476_i_0);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    \serCON_WRITE_PROC.sercon_8_0_0[3]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => \sercon[6]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => N_1064, D => N_189, Y => \sercon_8_0_0[3]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \fsmsync_ns_i_0[6]\ : CFG4
      generic map(INIT => x"5C5F")

      port map(A => \SDAInt\, B => \COREI2C_0_4_INT[0]\, C => 
        \fsmsync[1]_net_1\, D => \sercon[4]_net_1\, Y => 
        \fsmsync_ns_i_0[6]_net_1\);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[26]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_18_s5_1_0, Y => 
        \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \CLK_COUNTER1_PROC.un1_bclke_1.CO2\ : CFG3
      generic map(INIT => x"01")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[21]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \sersta_RNI25TS1[3]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        seradr0apb(6), Y => N_1220);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_3_601_0_1, D => N_1717, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_ns_0_a4[5]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => \pedetect\, B => \SCLSCL\, C => un115_fsmdet, 
        D => \fsmmod[1]_net_1\, Y => N_1058);
    
    \fsmmod_ns_0_a4[0]\ : CFG4
      generic map(INIT => x"AAA2")

      port map(A => \fsmmod[6]_net_1\, B => \starto_en\, C => 
        N_1040, D => N_64, Y => N_1048);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \COREI2C_0_4_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \ack\, B => N_2177, C => N_133, D => 
        fsmsta_8_28_307_a3_0_1, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \sersta_32_i_a2_7[3]\, D => \COREI2C_0_4_INT[0]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    un1_fsmsta_1_i_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        Y => \un1_fsmsta_1_i_0_o2_0\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"0B00")

      port map(A => bclke, B => \PCLK_count1_ov_1_sqmuxa_1\, C
         => \un1_PCLK_count1_0_sqmuxa\, D => PCLK_count2_ov_6_1, 
        Y => \PCLK_count1_1_sqmuxa\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \ack\, B => \fsmsta[23]_net_1\, C => 
        \adrcompen\, D => \adrcomp\, Y => fsmsta_8_5_555_a3_0_1);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_4_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        PCLK_count2_ov_6_1, C => CO1, D => \PCLK_count1_1_sqmuxa\, 
        Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[16]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_1[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => un91_ens1, B => \sercon[6]_net_1\, C => 
        N_2179, Y => N_162);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        \un1_serdat_2_sqmuxa_1\, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    SCLO_int_RNIBS4D : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_4_SCLO[0]\, Y => 
        COREI2C_0_4_SCLO_i(0));
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[12]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => N_2186, B => N_2177, C => un136_framesync, D
         => N_82, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_863_i_0);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \sersta_32_4[1]\, B => m7_4, C => 
        \sersta_32_5[1]\, D => m7_5, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    un151_framesync_RNIAKC61 : CFG3
      generic map(INIT => x"DC")

      port map(A => \un151_framesync\, B => N_2177, C => N_191, Y
         => un1_fsmsta_10_i_0);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \fsmsync_ns_i_o3_0_i_o2[5]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_64, B => \fsmsync[5]_net_1\, Y => N_68);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[27]\, B => un136_framesync, C
         => N_2177, D => fsmsta_nxt_1_sqmuxa_24_s4_1_0, Y => 
        \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_bm[3]\ : CFG3
      generic map(INIT => x"6C")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[3]_net_1\, C => CO1_1, Y => 
        \framesync_7_enl_bm_0[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG4
      generic map(INIT => x"F0F4")

      port map(A => N_2177, B => fsmsta_8_5_555_a3_0_1, C => 
        N_1680, D => N_2181, Y => N_1665);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_4_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_4_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"7075")

      port map(A => \ack\, B => un13_adrcompen, C => 
        \adrcomp_2_sqmuxa_i_a2_1_5\, D => N_133, Y => N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_4_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_1\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[9]_net_1\, C
         => \adrcomp_2_sqmuxa_i_o2_1_1\, D => un135_ens1_3, Y => 
        un135_ens1_1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => N_1470);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_172, B => N_2177, C => fsmsta_8_5_555_a3_0, 
        D => N_1622_2, Y => N_1680);
    
    \fsmsta_RNO[19]\ : CFG4
      generic map(INIT => x"000B")

      port map(A => N_191, B => \fsmsta_8_i_a3_0[19]\, C => 
        N_2199, D => un136_framesync, Y => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \un151_framesync\, Y => 
        \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \COREI2C_0_4_INT[0]\, B => \sercon[5]_net_1\, 
        C => N_1041, D => \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => 
        N_1054);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_0\ : CFG4
      generic map(INIT => x"CFEE")

      port map(A => N_2182, B => N_2181, C => \fsmsta[9]_net_1\, 
        D => N_2177, Y => fsmsta_8_4_577_i_0);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[12]_net_1\, 
        C => \fsmsta[22]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        un25_fsmsta_1);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFBA")

      port map(A => un16_fsmmod, B => N_2177, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_RNIM9M01\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \nedetect\, B => \COREI2C_0_4_INT[0]\, C => 
        un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sn_N_10_mux);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_4_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO0, B => framesync_7_e2, C => 
        \framesync[1]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[1]\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F202")

      port map(A => \sercon_8_2[4]\, B => \fsmsta_cnst[0]\, C => 
        un5_penable, D => CoreAPB3_0_APBmslave0_PWDATA(4), Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[11]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => N_76, D => \fsmsync[4]_net_1\, Y => N_55_i_0);
    
    \FSMSTA_SYNC_PROC.un133_framesync\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \adrcomp\, B => \adrcompen\, C => un91_ens1, 
        D => \fsmsta[23]_net_1\, Y => un133_framesync);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un133_framesync, B => N_2181, Y => 
        un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \un1_PCLK_count1_0_sqmuxa\, D
         => \PCLK_count1_1_sqmuxa\, Y => \PCLK_count1_10[0]\);
    
    \serSTA_WRITE_PROC.sersta_32_4[0]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => \COREI2C_0_4_INT[0]\, B => N_127, C => 
        \fsmsta[9]_net_1\, Y => \sersta_32_4[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, Y => 
        un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO\ : CFG4
      generic map(INIT => x"C010")

      port map(A => \nedetect\, B => \COREI2C_0_4_INT[0]\, C => 
        bsd7_i_m_0, D => un105_ens1, Y => bsd7_i_m);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    un1_PCLK_count1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"CECC")

      port map(A => bclke, B => \PCLK_count1_0_sqmuxa_3\, C => 
        \PCLK_count1[3]_net_1\, D => CO2, Y => 
        \un1_PCLK_count1_0_sqmuxa_1\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => mst, B => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[0]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_enl_am_0[0]\);
    
    \fsmmod_ns_0_a4[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \nedetect\, B => un115_fsmdet, C => 
        \fsmmod[5]_net_1\, Y => N_1050);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    \un2_framesync_1_1.CO0\ : CFG3
      generic map(INIT => x"C8")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        un70_fsmsta, Y => CO0);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"22EF")

      port map(A => \COREI2C_0_4_SDAO[0]\, B => N_2177, C => 
        \fsmsta[22]_net_1\, D => \fsmsta[20]_net_1\, Y => 
        fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0045")

      port map(A => N_1064, B => \fsmmod[2]_net_1\, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \un5_penable_2\, B => N_8_0, C => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), D => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    un1_PCLK_count1_0_sqmuxa_1_0 : CFG4
      generic map(INIT => x"080C")

      port map(A => \sercon[0]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => CO2, D => ANC2, Y => 
        \un1_PCLK_count1_0_sqmuxa_1_0\);
    
    \sersta_RNIMOSS1[0]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1[3]\, C => \sersta[0]_net_1\, D => 
        \COREI2C_0_4_INT[0]\, Y => N_1217);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \sersta_RNIU0TS1[2]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        seradr0apb(5), Y => N_1219);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => \sercon[5]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    \serCON_WRITE_PROC.un5_penable_2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CONFIG_rega20_2, B => 
        CoreAPB3_0_APBmslave0_PADDR(1), C => un3_penable_1, D => 
        un105_ens1_3, Y => \un5_penable_2\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"4440")

      port map(A => un16_fsmmod, B => PCLK_count2_ov_6_0_a2_1_3, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    un1_counter_rst_3 : CFG2
      generic map(INIT => x"B")

      port map(A => \PCLK_count1_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, Y => \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_4_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"ACAA")

      port map(A => \fsmsta[13]_net_1\, B => 
        \COREI2C_0_4_SDAO[0]\, C => N_2177, D => N_2196, Y => 
        N_82);
    
    \fsmsta_RNO[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1656, B => N_2186, C => N_2181, D => N_124, 
        Y => N_1774_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_4_SDAO[0]\, Y => 
        N_172);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_m1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        \serdat_0_sqmuxa\, Y => bsd7_tmp_6_m1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_4, B => N_145_2, C => 
        N_2177, D => fsmsta_8_20_379_i_0_a3_5, Y => N_145);
    
    adrcomp : SLE
      port map(D => N_2176, CLK => FAB_CCC_GL0, EN => 
        adrcomp_2_sqmuxa_i_0_3, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[19]_net_1\, 
        C => \fsmsta[4]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_4);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \fsmmod[0]_net_1\, B => \fsmdet[3]_net_1\, C
         => \fsmdet[1]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        N_1717);
    
    un1_fsmsta_i_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[18]_net_1\, 
        Y => un135_ens1_7);
    
    \serCON_WRITE_PROC.un91_ens1_0_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2177, B => \pedetect\, Y => un91_ens1);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0_RNIPO2K\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[20]_net_1\, 
        C => un57_fsmsta_1_0, Y => N_191);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[10]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[9]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \PCLKint\, B => \PCLKint_ff\, C => N_1586_1, 
        D => \fsmmod[2]_net_1\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \COREI2C_0_4_INT[0]\, B => N_1041, C => 
        \sercon[4]_net_1\, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[26]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, Y
         => N_145_2);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \sersta_RNI69TS1[4]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        seradr0apb(7), Y => N_1221);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => N_1665, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_68, B => \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1050, Y => \fsmmod_ns[1]\);
    
    \serdat_RNI4TB11[4]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(4), B => \serdat[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1[4]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_4_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    mst_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, Y
         => mst);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => un135_ens1_2, C => 
        \un151_framesync\, D => un57_fsmsta_1_0, Y => un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_2181, B => fsmsta_8_2_647_i_0_0, C => 
        N_1656, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_3\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[16]_net_1\, C
         => \fsmsta[20]_net_1\, D => \fsmsta[8]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    un1_PCLK_count1_0_sqmuxa : CFG4
      generic map(INIT => x"EEEF")

      port map(A => \un1_PCLK_count1_0_sqmuxa_1\, B => 
        \un1_PCLK_count1_0_sqmuxa_0\, C => \sercon[7]_net_1\, D
         => \un1_PCLK_count1_0_sqmuxa_1_0\, Y => 
        \un1_PCLK_count1_0_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => un1_fsmsta_10_i_0, B => \fsmsta[22]_net_1\, C
         => un136_framesync, D => \fsmsta_nxt_9_m[22]\, Y => 
        \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_3, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \framesync_7_enl_bm_0[0]\, B => 
        \framesync_7_enl_am_0[0]\, C => framesync_7_e2, Y => 
        \framesync_7[0]\);
    
    \sersta_RNIQSSS1[1]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1[4]\, C => \sersta[1]_net_1\, D => 
        \sercon[4]_net_1\, Y => N_1218);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_counter_rst_3\, D => 
        \un1_PCLK_count1_0_sqmuxa\, Y => \PCLK_count1_10[1]\);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG4
      generic map(INIT => x"F1F0")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_64, D => N_1002_3, Y => N_70);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        fsmsta_8_10_476_i_a6_1);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \bsd7_tmp\, B => \SCLInt\, C => 
        \COREI2C_0_4_INT[0]\, D => un57_fsmsta, Y => 
        bsd7_tmp_i_m_2);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"F0F8")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat_2_sqmuxa_1_0\, Y => 
        un1_serdat_2_sqmuxa_3);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \COREI2C_0_4_INT[0]\, B => N_1002, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_4_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.un25_framesync\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \sercon[5]_net_1\, B => \sercon[4]_net_1\, C
         => \COREI2C_0_4_INT[0]\, D => \un151_framesync\, Y => 
        un25_framesync);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"0C08")

      port map(A => un92_fsmsta, B => \pedetect\, C => un105_ens1, 
        D => \un1_serdat40\, Y => \un1_serdat_2_sqmuxa_1\);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[10]_net_1\, C => 
        N_1657_2, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_172, B => N_2182, C => N_2193, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_1002_3, B => 
        \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[2]_net_1\, Y => N_1002);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[27]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_24_s4_1_0);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"0013")

      port map(A => N_1624, B => fsmsta_8_10_476_i_0, C => 
        fsmsta_8_10_476_i_a6_1, D => N_1622_2, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[3]_net_1\, B => \serdat[2]_net_1\, C
         => \serdat[1]_net_1\, D => \serdat[0]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta[11]_net_1\, C
         => \fsmsta[7]_net_1\, D => \fsmsta[23]_net_1\, Y => m7_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_172, B => \fsmsta[26]_net_1\, Y => 
        fsmsta_nxt_1_sqmuxa_18_s5_1_0);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_4_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \serdat_RNIHLIV[5]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[5]_net_1\, B => \sercon[5]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3430")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1586_1, D => un1_fsmmod, Y => N_1624);
    
    adrcomp_2_sqmuxa_i_o2 : CFG2
      generic map(INIT => x"D")

      port map(A => mst, B => \fsmsta[23]_net_1\, Y => N_95);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_4_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        \COREI2C_0_4_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_1054, B => N_1046, C => 
        \fsmmod_ns_i_0[2]_net_1\, D => un115_fsmdet, Y => 
        N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \CLK_COUNTER1_PROC.un12_pclk_count1_1.CO3\ : CFG4
      generic map(INIT => x"777F")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => un12_pclk_count1);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    SDAO_int_RNI1B4 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_4_SDAO[0]\, Y => 
        COREI2C_0_4_SDAO_i(0));
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_1[3]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => un74_ens1, B => \adrcomp\, C => N_162, D => 
        N_163_2, Y => \sercon_8_0_1[3]\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[23]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_5);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNIVGE41 : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        \pedetect\, C => un136_framesync, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \serdat_RNIJNIV[6]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[6]_net_1\, B => \sercon[6]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_4_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => \PCLKint_ff\, D => \PCLKint\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => SDAO_int_7_0_275, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_4_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[19]_net_1\, 
        C => \fsmsta[20]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_2181, B => N_145, C => 
        fsmsta_8_20_379_i_0_o2_0, D => N_166, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_sm0, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[15]_net_1\, C
         => \fsmsta[17]_net_1\, D => \fsmsta[6]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    PCLKint_ff_RNILFDD : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \fsmsync_ns_i_a3_1_0_a2_1[2]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[0]_net_1\, Y
         => \fsmsync_ns_i_a3_1_0_a2_1[2]_net_1\);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_9_509_0_1, D => N_1717, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => N_126, B => N_2181, C => un133_framesync, D
         => N_80, Y => N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"FBF8")

      port map(A => \PWDATA_i_m_1[7]\, B => un105_ens1, C => 
        \fsmdet[3]_net_1\, D => bsd7_tmp_i_m_2, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \PCLKint\, B => \un151_framesync\, C => 
        \PCLKint_ff\, Y => \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[4]_net_1\, C => N_1657_2, 
        D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"5444")

      port map(A => un115_fsmdet, B => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, C => \fsmmod[3]_net_1\, D
         => N_1034, Y => \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FDFF")

      port map(A => m7_4, B => \sersta_32_3[0]\, C => 
        \sersta_32_4[0]\, D => m7_5, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => un135_ens1_1, C
         => un135_ens1_7, D => un135_ens1_2, Y => un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        un1_serdat_2_sqmuxa_3, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0301")

      port map(A => \fsmmod[6]_net_1\, B => \fsmmod[2]_net_1\, C
         => \fsmmod[0]_net_1\, D => \adrcomp\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    un1_serdat_2_sqmuxa_1_0 : CFG4
      generic map(INIT => x"00EF")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => un57_fsmsta, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1_0\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => \bsd7_tmp\, B => bsd7_tmp_6_m1, C => 
        bsd7_tmp_6_sm0, D => bsd7_tmp_6_sn_N_10_mux, Y => 
        bsd7_tmp_6);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un3_penable_1, B => N_43, C => un105_ens1_0, 
        D => un105_ens1_3, Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_4_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \fsmsync_RNO[1]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_1007, B => \fsmsync_ns_i_0[6]_net_1\, C => 
        N_1002, Y => N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1058, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \fsmsta[12]_net_1\, B => \COREI2C_0_4_INT[0]\, 
        C => \fsmsta[28]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_4_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_am[3]\ : CFG4
      generic map(INIT => x"FF07")

      port map(A => un70_fsmsta, B => un19_framesync, C => 
        un25_framesync, D => framesync_7_sm0, Y => 
        \framesync_7_enl_am_0[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[5]_net_1\, B => \fsmsync[2]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG4
      generic map(INIT => x"0307")

      port map(A => \fsmmod[0]_net_1\, B => \nedetect\, C => 
        \fsmmod[4]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \fsmmod_ns_i_0[2]_net_1\);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_2181, B => \ack\, C => un13_adrcompen, Y
         => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_3);
    
    adrcomp_2_sqmuxa_i_o2_1_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, Y
         => \adrcomp_2_sqmuxa_i_o2_1_1\);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_3 is

    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0);
          COREI2C_0_4_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 1);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 13);
          MSS_READY                                  : in    std_logic;
          FAB_CCC_GL0                                : in    std_logic;
          un3_penable                                : in    std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          BIBUF_COREI2C_0_4_SDA_IO_Y                 : in    std_logic;
          BIBUF_COREI2C_0_4_SCL_IO_Y                 : in    std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic;
          un3_penable_1                              : in    std_logic;
          un105_ens1_3                               : in    std_logic;
          un5_penable_2                              : out   std_logic;
          bclke                                      : in    std_logic;
          N_8_0                                      : in    std_logic;
          N_43                                       : in    std_logic;
          un105_ens1_0                               : in    std_logic
        );

end COREI2C_3;

architecture DEF_ARCH of COREI2C_3 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_3
    port( COREI2C_0_4_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_INT                            : out   std_logic_vector(0 to 0);
          seradr0apb                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 1) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 13) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          BIBUF_COREI2C_0_4_SDA_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_4_SCL_IO_Y                 : in    std_logic := 'U';
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic := 'U';
          un3_penable_1                              : in    std_logic := 'U';
          un105_ens1_3                               : in    std_logic := 'U';
          un5_penable_2                              : out   std_logic;
          bclke                                      : in    std_logic := 'U';
          N_8_0                                      : in    std_logic := 'U';
          N_43                                       : in    std_logic := 'U';
          un105_ens1_0                               : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_3
	Use entity work.COREI2CREAL_6_3(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_3
      port map(COREI2C_0_4_SDAO_i(0) => COREI2C_0_4_SDAO_i(0), 
        COREI2C_0_4_SCLO_i(0) => COREI2C_0_4_SCLO_i(0), 
        COREI2C_0_4_INT(0) => COREI2C_0_4_INT(0), seradr0apb(7)
         => \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14), 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13), 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, N_1218 => N_1218, N_1219 => 
        N_1219, N_1217 => N_1217, N_1220 => N_1220, N_1221 => 
        N_1221, BIBUF_COREI2C_0_4_SDA_IO_Y => 
        BIBUF_COREI2C_0_4_SDA_IO_Y, BIBUF_COREI2C_0_4_SCL_IO_Y
         => BIBUF_COREI2C_0_4_SCL_IO_Y, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, CONFIG_rega20_2 => 
        CONFIG_rega20_2, un3_penable_1 => un3_penable_1, 
        un105_ens1_3 => un105_ens1_3, un5_penable_2 => 
        un5_penable_2, bclke => bclke, N_8_0 => N_8_0, N_43 => 
        N_43, un105_ens1_0 => un105_ens1_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2CREAL_6_1 is

    port( COREI2C_0_2_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          seradr0apb                   : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          bclke                        : in    std_logic;
          N_1218                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_2_SCL_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_2_SDA_IO_Y   : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un3_penable_1                : in    std_logic;
          un105_ens1_1                 : in    std_logic;
          N_40                         : in    std_logic;
          un5_penable_1                : in    std_logic
        );

end COREI2CREAL_6_1;

architecture DEF_ARCH of COREI2CREAL_6_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREI2C_0_2_SDAO[0]\, \COREI2C_0_2_SCLO[0]\, 
        \SCLInt\, SCLInt_i_0, \fsmdet[3]_net_1\, \fsmdet_i_0[3]\, 
        \SCLI_ff_reg[0]_net_1\, GND_net_1, \SCLI_ff_reg_3[0]\, 
        VCC_net_1, \SCLI_ff_reg[1]_net_1\, \SCLI_ff_reg_3[1]\, 
        \SCLI_ff_reg[2]_net_1\, \SCLI_ff_reg_3[2]\, 
        \SDAI_ff_reg[0]_net_1\, \SDAI_ff_reg_4[0]\, 
        \SDAI_ff_reg[1]_net_1\, \SDAI_ff_reg_4[1]\, 
        \SDAI_ff_reg[2]_net_1\, \SDAI_ff_reg_4[2]\, 
        \indelay[0]_net_1\, N_57_i_0, \indelay[1]_net_1\, 
        N_55_i_0, \indelay[2]_net_1\, N_53_i_0, 
        \indelay[3]_net_1\, N_51_i_0, \PCLK_count2[0]_net_1\, 
        \PCLK_count2_3[0]\, \PCLK_count2[1]_net_1\, 
        \PCLK_count2_3[1]\, \PCLK_count2[2]_net_1\, 
        \PCLK_count2_3[2]\, \PCLK_count2[3]_net_1\, 
        \PCLK_count2_3[3]\, \framesync[0]_net_1\, 
        \framesync_7[0]\, \framesync[1]_net_1\, \framesync_7[1]\, 
        \framesync[2]_net_1\, \framesync_7[2]\, 
        \framesync[3]_net_1\, \framesync_7[3]\, \sercon[0]_net_1\, 
        un5_penable, \sercon[1]_net_1\, \sercon[2]_net_1\, 
        \COREI2C_0_2_INT[0]\, \sercon_9[3]\, \sercon[4]_net_1\, 
        \sercon_9[4]\, \sercon[5]_net_1\, \sercon[6]_net_1\, 
        \sercon[7]_net_1\, \PCLK_count1[0]_net_1\, 
        \PCLK_count1_10[0]\, \PCLK_count1[1]_net_1\, 
        \PCLK_count1_10[1]\, \PCLK_count1[2]_net_1\, 
        \PCLK_count1_10[2]\, \PCLK_count1[3]_net_1\, 
        \PCLK_count1_10[3]\, \serdat[2]_net_1\, \serdat_9[2]\, 
        \un1_serdat_2_sqmuxa_1\, \serdat[3]_net_1\, \serdat_9[3]\, 
        \serdat[4]_net_1\, \serdat_9[4]\, \serdat[5]_net_1\, 
        \serdat_9[5]\, \serdat[6]_net_1\, \serdat_9[6]\, 
        \serdat[7]_net_1\, \serdat_9[7]\, \serdat[0]_net_1\, 
        \serdat_9[0]\, \serdat[1]_net_1\, \serdat_9[1]\, 
        \sersta[0]_net_1\, \sersta_32[0]\, \sersta[1]_net_1\, 
        \sersta_32[1]\, \sersta[2]_net_1\, \sersta_32[2]\, 
        \sersta[3]_net_1\, N_99_i_0, \sersta[4]_net_1\, N_100_i_0, 
        \fsmsta[14]_net_1\, N_36_i_0, un1_ens1_pre_1_sqmuxa_i_0, 
        \fsmsta[13]_net_1\, N_34_i_0, \fsmsta[12]_net_1\, 
        N_1774_i_0, \fsmsta[11]_net_1\, N_1751_i_0, 
        \fsmsta[10]_net_1\, N_1701, \fsmsta[9]_net_1\, N_2172_i_0, 
        \fsmsta[8]_net_1\, fsmsta_8_5_555_0, \fsmsta[7]_net_1\, 
        \fsmsta_8[7]\, \fsmsta[6]_net_1\, N_44_i_0, 
        \fsmsta[5]_net_1\, N_42_i_0, \fsmsta[4]_net_1\, N_1631, 
        \fsmsta[3]_net_1\, N_1622_i_0, \fsmsta[2]_net_1\, 
        N_1604_i_0, \fsmsta[1]_net_1\, N_1586_i_0, 
        \fsmsta[0]_net_1\, N_1549, \fsmsta[29]_net_1\, 
        \fsmsta_8[29]\, \fsmsta[28]_net_1\, \fsmsta_8[28]\, 
        \fsmsta[27]_net_1\, \fsmsta_8[27]\, \fsmsta[26]_net_1\, 
        \fsmsta_8[26]\, \fsmsta[25]_net_1\, N_2175_i_0, 
        \fsmsta[24]_net_1\, \fsmsta_8[24]\, \fsmsta[23]_net_1\, 
        N_1543_i_0, \fsmsta[22]_net_1\, \fsmsta_8[22]\, 
        \fsmsta[21]_net_1\, \fsmsta_8[21]\, \fsmsta[20]_net_1\, 
        N_1520_i_0, \fsmsta[19]_net_1\, N_2174_i_0, 
        \fsmsta[18]_net_1\, \fsmsta_8[18]\, \fsmsta[17]_net_1\, 
        N_2173_i_0, \fsmsta[16]_net_1\, \fsmsta_8[16]\, 
        \fsmsta[15]_net_1\, N_1470, \ack\, ack_7, N_1449, 
        SDAO_int_1_sqmuxa_i_0, \bsd7_tmp\, bsd7_tmp_6, \bsd7\, 
        bsd7_9_iv_i_0, \adrcomp\, N_2176_i_0, 
        adrcomp_2_sqmuxa_i_0_1, \PCLKint\, PCLKint_3, 
        un1_pclkint4_i_0, \ack_bit\, \ack_bit_1_sqmuxa\, 
        \busfree\, un105_fsmdet, \adrcompen\, 
        \adrcompen_0_sqmuxa\, adrcompen_2_sqmuxa_i_0, \SCLSCL\, 
        \fsmmod[1]_net_1\, SCLSCL_1_sqmuxa_i_0, \SDAInt\, 
        un1_rtn_4_1, un1_rtn_3_1, \nedetect\, \nedetect_0_sqmuxa\, 
        rtn_i_0, \pedetect\, \pedetect_0_sqmuxa\, rtn_1, 
        \starto_en\, N_40_i_0, N_60, \fsmdet[0]_net_1\, N_867_i_0, 
        \fsmsync[7]_net_1\, \fsmsync_ns[0]\, \fsmsync[6]_net_1\, 
        N_966_i_0, \fsmsync[5]_net_1\, N_968_i_0, 
        \fsmsync[4]_net_1\, N_970_i_0, \fsmsync[3]_net_1\, 
        N_972_i_0, \fsmsync[2]_net_1\, N_974_i_0, 
        \fsmsync[1]_net_1\, N_976_i_0, \fsmdet[6]_net_1\, 
        \fsmdet[5]_net_1\, N_857_i_0, \fsmdet[4]_net_1\, 
        N_859_i_0, N_861_i_0, \fsmdet[2]_net_1\, N_863_i_0, 
        \fsmdet[1]_net_1\, N_865_i_0, \fsmmod[6]_net_1\, 
        \fsmmod_ns[0]\, \fsmmod[5]_net_1\, \fsmmod_ns[1]\, 
        \fsmmod[4]_net_1\, N_1026_i_0, \fsmmod[3]_net_1\, 
        \fsmmod_ns[3]\, \fsmmod[2]_net_1\, N_1029_i_0, 
        \fsmmod_ns[5]\, \fsmmod[0]_net_1\, N_1032_i_0, 
        un149_ens1_i_0, \PCLKint_ff\, PCLKint_ff_2, 
        \PCLK_count1_ov\, \PCLK_count1_1_sqmuxa\, 
        \PCLK_count2_ov\, PCLK_count2_ov_6, PCLK_count2_ov_6_1, 
        \un1_PCLK_count1_0_sqmuxa\, CO1, un13_adrcompen, 
        \adrcomp_2_sqmuxa_i_a2_1_5\, N_2187, un57_fsmsta, 
        \un1_serdat40\, \un1_serdat_2_sqmuxa_1_0\, N_66, N_84, 
        \sersta_32_5[2]\, un16_fsmmod, N_1586_1, N_2181, 
        un105_ens1, N_2177, N_2173_i_1, N_133, un1_fsmmod, 
        N_36_i_1, un136_framesync, N_2196, N_2186, 
        \fsmsta_8_1[24]\, un57_fsmsta_1_0, N_172, 
        \PCLK_count1_0_sqmuxa_4\, \PCLK_count1_0_sqmuxa_3\, 
        \un1_PCLK_count1_0_sqmuxa_0\, 
        \un1_PCLK_count1_0_sqmuxa_1_0\, CO2, \fsmsta_cnst[0]\, 
        fsmsta_8_9_509_0_1, N_1717, fsmsta_8_9_509_0, N_1658_1, 
        N_1652, fsmsta_8_3_601_0_1, fsmsta_8_3_601_0, 
        \un1_pclk_count1_ov_1_1\, \un1_pclk_count1_ov_1\, 
        \PRDATA_3_1_1[4]\, \PRDATA_3_1_1[7]\, \PRDATA_3_1_1[3]\, 
        \PRDATA_3_1_1[5]\, \PRDATA_3_1_1[6]\, \fsmsta_8_ns_1[29]\, 
        \fsmsta_8_ns_1[28]\, \fsmsta_8_ns_1[16]\, un133_framesync, 
        \fsmsta_8_ns_1[18]\, framesync_7_sm0, 
        \framesync_7_enl_ns_1[3]\, \framesync_7_m0[3]\, 
        framesync_7_e2, CO0, N_2179, N_161_2, un70_fsmsta, 
        fsmsta_8_10_476_i_a6_0, PCLK_count2_ov_6_0_a2_1_0, 
        \fsmsta_nxt_9_m_0[27]\, \fsmsta_nxt_9_m_0[26]\, 
        \sersta_32_2[0]\, un111_fsmdet_0, \sersta_32_i_a2_5[3]\, 
        un139_ens1_0, N_997, fsmsta_8_20_379_i_0_a3_3, 
        \un1_fsmsta_1_i_0_o2_0\, un26_adrcompen_6, un135_ens1_2, 
        N_67, N_64, N_153_1, N_23, N_127, mst, N_2178, N_1196, 
        N_1197, N_1198, SDAO_int_7_0_275_1, 
        \adrcomp_2_sqmuxa_i_a3_3\, SDAO_int_7_0_275_a5_0, 
        un141_ens1_2, \SDAO_int_1_sqmuxa_3\, 
        \adrcomp_2_sqmuxa_i_a2_1_2\, \adrcomp_2_sqmuxa_i_a2_1_0\, 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\, fsmsta_8_5_555_a3_0_1, 
        fsmsta_8_5_555_a3_0, \sersta_32_3[0]\, \sersta_32_5[1]\, 
        \sersta_32_4[1]\, \fsmmod_ns_i_a4_1_0[2]_net_1\, 
        fsmsta_8_20_379_i_0_a3_4, fsmsta_8_20_379_i_0_a3_3_0, 
        \sersta_32_i_a2_7[4]\, \sersta_32_i_a2_6[4]\, 
        \sersta_32_4[2]\, un135_ens1_5, un135_ens1_4, 
        un135_ens1_3, un57_fsmsta_0, un25_fsmsta_2, 
        \sersta_32_i_a2_8[3]\, \sersta_32_i_a2_7[3]\, 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, 
        \adrcomp_2_sqmuxa_i_o2_1_3\, m7_3, un13_adrcompen_4, 
        \PCLK_count1_ov_1_sqmuxa_1\, un19_framesync_1, 
        \PCLK_count1_0_sqmuxa_1_1\, N_1064, un12_pclk_count1, 
        un33_fsmsta, PCLK_count2_ov_6_0_a2_1_4_tz, N_76, CO2_0, 
        \un1_pclk_count1_ov\, CO1_0, N_1040, N_117_1, N_1049, 
        N_1034, un149_framesync, N_2182, 
        \adrcomp_2_sqmuxa_i_a3_4\, \fsmmod_ns_i_0[2]_net_1\, 
        \SDAO_int_1_sqmuxa_4\, \adrcomp_2_sqmuxa_i_a2_1_4\, 
        PCLK_count2_ov_6_0_a2_1_3, \adrcomp_2_sqmuxa_i_0_0_0\, 
        \sercon_8_0_a3_1_0[3]\, \sersta_32_i_a2_9[4]\, 
        \sercon_8_2[4]\, \sersta_32_7[2]\, \sersta_32_i_a2_10[3]\, 
        N_72_mux, un25_fsmsta, N_1002, 
        fsmsta_nxt_1_sqmuxa_18_s5_1, N_104, N_2192, 
        fsmsta_nxt_1_sqmuxa_24_s4_1, \fsmsta_8_0_a2_1[7]\, N_134, 
        N_1041, N_1622_2, un74_ens1, N_63, \un1_pclk_count191\, 
        N_995, N_130, N_1732, N_1656, N_2171, \un1_fsmsta_6\, 
        N_2193, N_120, N_124, fsmsta_8_10_476_i_1, 
        fsmsta_8_28_307_a3_0_1, \SDAO_int_1_sqmuxa_7\, 
        \fsmsync_ns_i_1[6]_net_1\, N_163, un135_ens1, N_165, 
        N_1054, N_157, un115_fsmdet, \framesync_1_sqmuxa\, 
        \fsmsta_nxt_9_m[21]\, \fsmsta_nxt_9_m[22]\, 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, N_1046, N_70, N_1048, 
        N_126, N_1657_2, N_1624, \framesync_0_sqmuxa\, N_1060, 
        N_193, \fsmsta_8_i_0[25]\, fsmsta_8_4_577_i_0, N_82, N_80, 
        bsd7_i_m_0, bsd7_tmp_i_m_2, fsmsta_8_20_379_i_0_o2_0, 
        \sercon_8_0_1[3]\, \fsmsync_ns_0_0_1[0]_net_1\, 
        fsmsta_8_23_351_i_0_1, \un1_ens1_pre_1_sqmuxa_0_a2_1\, 
        N_1680, N_145, N_1058, N_1050, N_1465, N_166, 
        \fsmsync_ns_i_0_1_tz[3]_net_1\, N_86, N_1059_1, 
        un1_fsmsta_10_i_0, un92_fsmsta, N_2199, \PWDATA_i_m_1[7]\, 
        \sercon_8_0_2[3]\, fsmsta_8_2_647_i_0_0, N_1486, N_161, 
        CO1_1, \framesync_7_m2[3]\, \serdat_0_sqmuxa\, 
        un134_fsmsta, N_1466, bsd7_tmp_6_sn_N_10_mux, N_152, 
        bsd7_tmp_6_m1, bsd7_tmp_6_sm0, \un1_counter_rst_3\, 
        bsd7_9_iv_1, bsd7_i_m, un1_serdat_2_sqmuxa_1_1
         : std_logic;

begin 

    COREI2C_0_2_INT(0) <= \COREI2C_0_2_INT[0]\;

    \SDAO_INT_WRITE_PROC.un33_fsmsta_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un33_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[21]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_193, B => N_2177, Y => un1_fsmsta_10_i_0);
    
    \sersta_RNO[3]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_23, B => \sersta_32_i_a2_5[3]\, C => 
        \sersta_32_i_a2_10[3]\, D => \sersta_32_i_a2_8[3]\, Y => 
        N_99_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2171, B => \sercon[2]_net_1\, Y => N_126);
    
    \FSMMOD_SYNC_PROC.un115_fsmdet\ : CFG4
      generic map(INIT => x"BBFB")

      port map(A => \fsmdet[1]_net_1\, B => \sercon[6]_net_1\, C
         => un111_fsmdet_0, D => N_2177, Y => un115_fsmdet);
    
    \sercon[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[1]_net_1\);
    
    \fsmmod_ns_0_o3_1[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \PCLKint\, B => \PCLKint_ff\, Y => N_64);
    
    adrcomp_2_sqmuxa_i_a2_1_5 : CFG4
      generic map(INIT => x"9000")

      port map(A => \serdat[0]_net_1\, B => seradr0apb(1), C => 
        \adrcomp_2_sqmuxa_i_a2_1_4\, D => 
        \adrcomp_2_sqmuxa_i_a2_1_0\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_5\);
    
    un1_fsmsta_nxt_0_sqmuxa_i : CFG3
      generic map(INIT => x"BA")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_153_1, 
        Y => N_2171);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7_3\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[27]_net_1\, 
        C => \fsmsta[4]_net_1\, D => \fsmsta[15]_net_1\, Y => 
        m7_3);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_1\ : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmsta[23]_net_1\, B => un1_fsmmod, C => 
        N_193, Y => N_166);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns[3]\ : CFG4
      generic map(INIT => x"CCFA")

      port map(A => framesync_7_sm0, B => 
        \framesync_7_enl_ns_1[3]\, C => \framesync_7_m0[3]\, D
         => framesync_7_e2, Y => \framesync_7[3]\);
    
    \fsmdet[1]\ : SLE
      port map(D => N_865_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[1]_net_1\);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet_3_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \fsmmod[2]_net_1\, B => \SCLInt\, C => N_64, 
        Y => N_1064);
    
    adrcomp_2_sqmuxa_i_a2_1_4 : CFG4
      generic map(INIT => x"0090")

      port map(A => \serdat[3]_net_1\, B => seradr0apb(4), C => 
        \adrcomp_2_sqmuxa_i_a2_1_2\, D => un26_adrcompen_6, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_4\);
    
    SDAInt : SLE
      port map(D => \SDAI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_4_1, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SDAInt\);
    
    starto_en : SLE
      port map(D => N_40_i_0, CLK => FAB_CCC_GL0, EN => N_60, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \starto_en\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \bsd7\, Y => bsd7_i_m_0);
    
    \fsmsync_ns_0_0_a2_2_1[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmmod[4]_net_1\, Y => N_117_1);
    
    \un1_PCLK_count2_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \PCLK_count2[1]_net_1\, C => \PCLK_count1_ov\, Y => CO1_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_a4_2\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_1656, B => \fsmdet[1]_net_1\, Y => N_1657_2);
    
    \serdat[4]\ : SLE
      port map(D => \serdat_9[4]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0[7]\ : CFG4
      generic map(INIT => x"3302")

      port map(A => N_126, B => un136_framesync, C => \SDAInt\, D
         => \fsmsta_8_0_a2_1[7]\, Y => \fsmsta_8[7]\);
    
    \fsmsta[4]\ : SLE
      port map(D => N_1631, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[4]_net_1\);
    
    \SCLI_ff_reg[1]\ : SLE
      port map(D => \SCLI_ff_reg_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[1]_net_1\);
    
    pedetect : SLE
      port map(D => \pedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pedetect\);
    
    \fsmmod[4]\ : SLE
      port map(D => N_1026_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[4]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[14]_net_1\, 
        C => un25_fsmsta_2, D => N_2178, Y => un25_fsmsta);
    
    \serSTA_WRITE_PROC.sersta_32[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \sersta_32_5[2]\, B => \sersta_32_7[2]\, C
         => un135_ens1_2, D => \un1_fsmsta_1_i_0_o2_0\, Y => 
        \sersta_32[2]\);
    
    \fsmmod_ns_0_a4_0_4[3]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1041, B => \fsmmod_ns_0_a4_0_4_2[3]_net_1\, 
        C => N_1040, Y => \fsmmod_ns_0_a4_0_4[3]_net_1\);
    
    un7_fsmsta_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[20]_net_1\, B => \fsmsta[22]_net_1\, 
        Y => N_2178);
    
    \fsmmod_ns_0[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_1064, B => N_1049, C => un115_fsmdet, D => 
        N_1048, Y => \fsmmod_ns[0]\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[1]_net_1\, Y
         => N_1586_1);
    
    adrcomp_2_sqmuxa_i_o2_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[23]_net_1\, B => 
        \adrcomp_2_sqmuxa_i_o2_1_3\, C => \fsmsta[3]_net_1\, D
         => \fsmsta[13]_net_1\, Y => N_2192);
    
    \PRDATA_3[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(1), C => N_1197, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1215);
    
    ack : SLE
      port map(D => ack_7, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \ack\);
    
    \fsmsta[3]\ : SLE
      port map(D => N_1622_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[3]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[1]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \PCLK_count2[1]_net_1\, B => \PCLK_count1_ov\, 
        C => \PCLK_count2[0]_net_1\, D => PCLK_count2_ov_6_1, Y
         => \PCLK_count2_3[1]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0_1\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => N_2181, C => 
        \adrcompen\, D => \adrcomp\, Y => fsmsta_8_28_307_a3_0_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => un1_fsmmod, B => SDAO_int_7_0_275_a5_0, C => 
        N_1466, D => SDAO_int_7_0_275_1, Y => N_1449);
    
    \serdat[2]\ : SLE
      port map(D => \serdat_9[2]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_1\ : CFG4
      generic map(INIT => x"FAF3")

      port map(A => N_1658_1, B => \fsmsta[3]_net_1\, C => 
        N_1622_2, D => N_1586_1, Y => fsmsta_8_10_476_i_1);
    
    un1_pclk_count1_ov_1 : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[1]_net_1\, C => \sercon[7]_net_1\, D => 
        \un1_pclk_count1_ov_1_1\, Y => \un1_pclk_count1_ov_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1586_1, B => un139_ens1_0, Y => 
        framesync_7_sm0);
    
    un7_fsmsta_i_0_o2_RNILPDU : CFG3
      generic map(INIT => x"01")

      port map(A => N_2178, B => un57_fsmsta_1_0, C => 
        \un1_fsmsta_6\, Y => N_193);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[29]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[5]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[29]\, Y => 
        \fsmsta_8[29]\);
    
    \fsmsta_RNO[9]\ : CFG4
      generic map(INIT => x"003A")

      port map(A => \ack\, B => N_172, C => N_2177, D => 
        fsmsta_8_4_577_i_0, Y => N_2172_i_0);
    
    \fsmmod_ns_0_a4_0[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \fsmmod[1]_net_1\, B => \SCLSCL\, C => 
        \pedetect\, Y => N_1049);
    
    un1_PCLK_count1_0_sqmuxa_0 : CFG4
      generic map(INIT => x"FF10")

      port map(A => \sercon[7]_net_1\, B => \sercon[1]_net_1\, C
         => un12_pclk_count1, D => \PCLK_count1_0_sqmuxa_1_1\, Y
         => \un1_PCLK_count1_0_sqmuxa_0\);
    
    \fsmsta_RNO[25]\ : CFG4
      generic map(INIT => x"0007")

      port map(A => N_172, B => N_2177, C => \fsmsta_8_i_0[25]\, 
        D => un136_framesync, Y => N_2175_i_0);
    
    \ADRCOMP_WRITE_PROC.un26_adrcompen_6\ : CFG2
      generic map(INIT => x"6")

      port map(A => \serdat[6]_net_1\, B => seradr0apb(7), Y => 
        un26_adrcompen_6);
    
    adrcomp_2_sqmuxa_i_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        \framesync[2]_net_1\, D => \framesync[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a3_3\);
    
    \fsmsta[23]\ : SLE
      port map(D => N_1543_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[23]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[29]_net_1\, 
        C => \fsmsta[21]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_3[0]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_2[3]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \sercon[6]_net_1\, B => \adrcomp\, C => 
        N_1586_1, D => un74_ens1, Y => N_163);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_o4\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1652, D => un1_fsmmod, Y => N_1656);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0_1\ : CFG3
      generic map(INIT => x"4E")

      port map(A => \framesync[3]_net_1\, B => N_1652, C => 
        \framesync[0]_net_1\, Y => fsmsta_8_3_601_0_1);
    
    \fsmsta[7]\ : SLE
      port map(D => \fsmsta_8[7]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[7]_net_1\);
    
    \serdat_RNI2PF21[5]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(5), B => \serdat[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[5]\);
    
    \fsmsta_RNO_0[17]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \fsmsta[23]_net_1\, B => \ack\, C => N_133, D
         => un1_fsmmod, Y => N_2173_i_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_1\ : CFG4
      generic map(INIT => x"F7F3")

      port map(A => \adrcomp\, B => \sercon[6]_net_1\, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[6]_net_1\, Y => 
        SDAO_int_7_0_275_1);
    
    \serCON_WRITE_PROC.sercon_8_0_o2[3]\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmdet[3]_net_1\, D => N_1064, Y => N_134);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_2_SDA_IO_Y, Y => \SDAI_ff_reg_4[0]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2_0[3]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \indelay[0]_net_1\, B => \indelay[2]_net_1\, 
        Y => N_67);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        N_161_2, Y => N_161);
    
    SDAO_int_1_sqmuxa_4 : CFG4
      generic map(INIT => x"0002")

      port map(A => \sercon[6]_net_1\, B => un1_fsmmod, C => 
        \fsmmod[3]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        \SDAO_int_1_sqmuxa_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1586_1, B => \fsmsta[8]_net_1\, Y => 
        fsmsta_8_5_555_a3_0);
    
    \un1_PCLK_count1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \un1_PCLK_count1_0_sqmuxa\, C => \PCLK_count1[1]_net_1\, 
        Y => CO1);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_66, B => \indelay[2]_net_1\, Y => N_76);
    
    \indelay_RNO[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => \indelay[0]_net_1\, B => \fsmsync[4]_net_1\, 
        C => N_76, Y => N_57_i_0);
    
    \serCON_WRITE_PROC.sercon_9[3]\ : CFG4
      generic map(INIT => x"FE32")

      port map(A => \sercon_8_0_2[3]\, B => un5_penable, C => 
        N_161, D => CoreAPB3_0_APBmslave0_PWDATA(3), Y => 
        \sercon_9[3]\);
    
    PCLK_count1_0_sqmuxa_4 : CFG4
      generic map(INIT => x"0004")

      port map(A => \sercon[7]_net_1\, B => CO2_0, C => 
        \sercon[1]_net_1\, D => \sercon[0]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_4\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[18]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[18]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[18]\, Y => 
        \fsmsta_8[18]\);
    
    \fsmmod[3]\ : SLE
      port map(D => \fsmmod_ns[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[3]_net_1\);
    
    \CLK_COUNTER1_PROC.un1_pclk_count1_1.CO2\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2_0);
    
    \PCLK_count2[3]\ : SLE
      port map(D => \PCLK_count2_3[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[3]_net_1\);
    
    un1_rtn_4 : CFG3
      generic map(INIT => x"81")

      port map(A => \SDAI_ff_reg[2]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, C => \SDAI_ff_reg[0]_net_1\, Y
         => un1_rtn_4_1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[21]\);
    
    \fsmsta[27]\ : SLE
      port map(D => \fsmsta_8[27]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[27]_net_1\);
    
    \fsmsta[6]\ : SLE
      port map(D => N_44_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[6]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_0_a2_1[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[7]_net_1\, C => N_172, Y
         => \fsmsta_8_0_a2_1[7]\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6s2\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sm0);
    
    \serdat[7]\ : SLE
      port map(D => \serdat_9[7]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[7]_net_1\);
    
    PCLK_count1_ov_1_sqmuxa_1 : CFG3
      generic map(INIT => x"80")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \PCLK_count1_ov_1_sqmuxa_1\);
    
    \sercon[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_o2_0_0\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => \fsmsta[23]_net_1\, B => N_172, C => N_2177, 
        D => N_165, Y => fsmsta_8_20_379_i_0_o2_0);
    
    \serCON_WRITE_PROC.sercon_8_2[4]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \sercon[4]_net_1\, B => \fsmdet[1]_net_1\, C
         => \sercon[6]_net_1\, D => mst, Y => \sercon_8_2[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[28]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[28]\);
    
    un1_serdat40 : CFG4
      generic map(INIT => x"0015")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => un25_fsmsta, D => un57_fsmsta, Y => \un1_serdat40\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1[24]\ : CFG4
      generic map(INIT => x"0F77")

      port map(A => \SDAInt\, B => un57_fsmsta_1_0, C => N_172, D
         => N_2177, Y => \fsmsta_8_1[24]\);
    
    adrcomp_2_sqmuxa_i_0 : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \COREI2C_0_2_INT[0]\, B => N_2192, C => 
        \adrcomp_2_sqmuxa_i_0_0_0\, D => N_152, Y => 
        adrcomp_2_sqmuxa_i_0_1);
    
    \un2_framesync_1_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync_1_sqmuxa\, C => \framesync[1]_net_1\, Y => 
        CO1_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_a5_0_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => \fsmmod[5]_net_1\, B => \fsmmod[0]_net_1\, C
         => \fsmmod[2]_net_1\, Y => SDAO_int_7_0_275_a5_0);
    
    SCLSCL : SLE
      port map(D => \fsmmod[1]_net_1\, CLK => FAB_CCC_GL0, EN => 
        SCLSCL_1_sqmuxa_i_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLSCL\);
    
    \fsmsta_RNO[20]\ : CFG3
      generic map(INIT => x"10")

      port map(A => fsmsta_8_23_351_i_0_1, B => N_2181, C => 
        N_1656, Y => N_1520_i_0);
    
    \serDAT_WRITE_PROC.serdat_9[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(1), B => 
        un105_ens1, C => \serdat[0]_net_1\, Y => \serdat_9[1]\);
    
    busfree_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \fsmdet[3]_net_1\, Y => \fsmdet_i_0[3]\);
    
    \SCLI_ff_reg[0]\ : SLE
      port map(D => \SCLI_ff_reg_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[0]_net_1\);
    
    \PRDATA_1[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[0]_net_1\, Y
         => N_1196);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0_1\ : CFG3
      generic map(INIT => x"32")

      port map(A => \framesync[3]_net_1\, B => N_1658_1, C => 
        N_1652, Y => fsmsta_8_9_509_0_1);
    
    \fsmsync_RNO[6]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \fsmsync[7]_net_1\, B => \SCLInt\, C => 
        N_1002, Y => N_966_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i\ : CFG4
      generic map(INIT => x"0045")

      port map(A => bsd7_9_iv_1, B => \serdat[7]_net_1\, C => 
        bsd7_tmp_6_sn_N_10_mux, D => bsd7_i_m, Y => bsd7_9_iv_i_0);
    
    \indelay_RNO[2]\ : CFG4
      generic map(INIT => x"6A00")

      port map(A => \indelay[2]_net_1\, B => \indelay[1]_net_1\, 
        C => \indelay[0]_net_1\, D => \fsmsync[4]_net_1\, Y => 
        N_53_i_0);
    
    \fsmsta[21]\ : SLE
      port map(D => \fsmsta_8[21]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[21]_net_1\);
    
    \fsmsta[16]\ : SLE
      port map(D => \fsmsta_8[16]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[16]_net_1\);
    
    \PRDATA_1[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \sercon[2]_net_1\, B => \serdat[2]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1198);
    
    \fsmmod_ns_i_a4[6]\ : CFG3
      generic map(INIT => x"31")

      port map(A => \fsmmod[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => N_1034, Y => N_1060);
    
    \serSTA_WRITE_PROC.sersta_32_5[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta[4]_net_1\, C
         => \fsmsta[24]_net_1\, D => \fsmsta[25]_net_1\, Y => 
        \sersta_32_5[2]\);
    
    adrcomp_2_sqmuxa_i_a2_1_0 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(3), B => seradr0apb(2), C => 
        \serdat[2]_net_1\, D => \serdat[1]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_0\);
    
    SDAO_int_1_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => un25_fsmsta, B => \SDAO_int_1_sqmuxa_7\, C
         => \SDAO_int_1_sqmuxa_3\, D => \SDAO_int_1_sqmuxa_4\, Y
         => SDAO_int_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_a3_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta_cnst[0]\, B => \fsmdet[3]_net_1\, Y
         => N_1732);
    
    PCLKint_RNO : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLK_count2_ov\, Y
         => un1_pclkint4_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_0_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, Y => fsmsta_8_10_476_i_a6_0);
    
    adrcomp_2_sqmuxa_i_a3 : CFG4
      generic map(INIT => x"D000")

      port map(A => mst, B => \fsmsta[23]_net_1\, C => N_2187, D
         => \adrcomp_2_sqmuxa_i_a3_4\, Y => N_152);
    
    un1_fsmsta_nxt_0_sqmuxa_i_a3_1 : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[8]_net_1\, Y
         => N_153_1);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_11_454_i_a6_2_0_0_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_fsmmod, B => \fsmsta[23]_net_1\, Y => 
        N_2182);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[2]\ : CFG4
      generic map(INIT => x"7D28")

      port map(A => framesync_7_e2, B => CO1_1, C => 
        \framesync[2]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_0\ : CFG4
      generic map(INIT => x"4577")

      port map(A => \fsmsta[11]_net_1\, B => N_2177, C => N_2186, 
        D => N_120, Y => fsmsta_8_2_647_i_0_0);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_6[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[1]_net_1\, C
         => \fsmsta[8]_net_1\, D => \fsmsta[7]_net_1\, Y => 
        \sersta_32_i_a2_6[4]\);
    
    SCLO_int_RNO : CFG4
      generic map(INIT => x"5777")

      port map(A => \sercon[6]_net_1\, B => un141_ens1_2, C => 
        un139_ens1_0, D => un135_ens1, Y => un149_ens1_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[28]\ : CFG4
      generic map(INIT => x"8F80")

      port map(A => \fsmdet[3]_net_1\, B => \fsmmod[0]_net_1\, C
         => un136_framesync, D => \fsmsta_8_ns_1[28]\, Y => 
        \fsmsta_8[28]\);
    
    \fsmsta_RNO[1]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[1]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1586_i_0);
    
    un1_pclk_count1_ov : CFG3
      generic map(INIT => x"13")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        \sercon[7]_net_1\, C => \PCLK_count2[1]_net_1\, Y => 
        \un1_pclk_count1_ov\);
    
    \PCLK_count2[0]\ : SLE
      port map(D => \PCLK_count2_3[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[0]_net_1\);
    
    \FSMMOD_SYNC_PROC.un111_fsmdet_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fsmsta[23]_net_1\, B => \pedetect\, Y => 
        un111_fsmdet_0);
    
    adrcomp_2_sqmuxa_i_0_0_0 : CFG2
      generic map(INIT => x"E")

      port map(A => un16_fsmmod, B => N_1586_1, Y => 
        \adrcomp_2_sqmuxa_i_0_0_0\);
    
    \sersta[0]\ : SLE
      port map(D => \sersta_32[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[0]_net_1\);
    
    \PCLK_count1[3]\ : SLE
      port map(D => \PCLK_count1_10[3]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[3]_net_1\);
    
    \indelay[2]\ : SLE
      port map(D => N_53_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[2]_net_1\);
    
    \fsmsync[2]\ : SLE
      port map(D => N_974_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_o2_0[19]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2177, B => N_2178, Y => N_2193);
    
    \fsmdet_RNO[5]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[5]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_857_i_0);
    
    \fsmsta[24]\ : SLE
      port map(D => \fsmsta_8[24]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[24]_net_1\);
    
    \framesync[3]\ : SLE
      port map(D => \framesync_7[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[3]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[29]_net_1\, C => N_172, 
        Y => \fsmsta_8_ns_1[29]\);
    
    \indelay_RNO[3]\ : CFG4
      generic map(INIT => x"A060")

      port map(A => \indelay[3]_net_1\, B => \indelay[1]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_67, Y => N_51_i_0);
    
    framesync_1_sqmuxa : CFG3
      generic map(INIT => x"20")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, Y
         => \framesync_1_sqmuxa\);
    
    \CLKINT_WRITE_PROC.PCLKint_ff_2\ : CFG2
      generic map(INIT => x"D")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_ff_2);
    
    \serdat_RNI4RF21[6]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(6), B => \serdat[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[6]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        BIBUF_COREI2C_0_2_SCL_IO_Y, Y => \SCLI_ff_reg_3[0]\);
    
    \fsmmod_ns_0_a4_0_1[1]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => \starto_en\, B => N_64, C => N_1040, D => 
        un115_fsmdet, Y => N_1059_1);
    
    \CLKINT_WRITE_PROC.PCLKint_3\ : CFG2
      generic map(INIT => x"7")

      port map(A => PCLK_count2_ov_6_1, B => \PCLKint\, Y => 
        PCLKint_3);
    
    un1_fsmsta_1_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_fsmsta_1_i_0_o2_0\, B => 
        \fsmsta[12]_net_1\, Y => N_2186);
    
    \fsmsta[15]\ : SLE
      port map(D => N_1470, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[15]_net_1\);
    
    un1_fsmsta_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[17]_net_1\, B => \fsmsta[14]_net_1\, 
        C => \fsmsta[18]_net_1\, Y => N_2196);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[8]_net_1\, Y
         => un135_ens1_2);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[0]\ : CFG4
      generic map(INIT => x"6F60")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync_1_sqmuxa\, C => framesync_7_e2, D => 
        \framesync_7_m2[3]\, Y => \framesync_7[0]\);
    
    PCLK_count1_ov : SLE
      port map(D => \PCLK_count1_1_sqmuxa\, CLK => FAB_CCC_GL0, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1_ov\);
    
    \indelay[1]\ : SLE
      port map(D => N_55_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[1]_net_1\);
    
    \fsmsta[22]\ : SLE
      port map(D => \fsmsta_8[22]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[22]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsync[3]_net_1\, B => \fsmsync[6]_net_1\, 
        Y => PCLK_count2_ov_6_0_a2_1_0);
    
    \FSMMOD_COMB_PROC.un149_framesync\ : CFG3
      generic map(INIT => x"02")

      port map(A => \sercon[5]_net_1\, B => \fsmsta[29]_net_1\, C
         => \fsmsta[28]_net_1\, Y => un149_framesync);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[3]\ : CFG4
      generic map(INIT => x"48C0")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[3]_net_1\, D => \PCLK_count2[2]_net_1\, Y
         => \PCLK_count2_3[3]\);
    
    \PRDATA_3[0]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(0), C => N_1196, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1214);
    
    \serdat[0]\ : SLE
      port map(D => \serdat_9[0]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[0]_net_1\);
    
    \fsmsta[10]\ : SLE
      port map(D => N_1701, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[10]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[26]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \un1_fsmsta_6\, B => un136_framesync, C => 
        \fsmsta_nxt_9_m_0[26]\, D => fsmsta_nxt_1_sqmuxa_18_s5_1, 
        Y => \fsmsta_8[26]\);
    
    \serCON_WRITE_PROC.un74_ens1\ : CFG4
      generic map(INIT => x"0009")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un74_ens1);
    
    \fsmmod_RNI8TEI2[0]\ : CFG4
      generic map(INIT => x"EEEC")

      port map(A => \fsmdet[3]_net_1\, B => \fsmsta_cnst[0]\, C
         => \fsmmod[5]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        N_1622_2);
    
    \CLK_COUNTER1_PROC.un1_bclke_1.CO2\ : CFG3
      generic map(INIT => x"01")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \PCLK_count1[0]_net_1\, Y
         => CO2);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[21]\ : CFG4
      generic map(INIT => x"5540")

      port map(A => un136_framesync, B => un1_fsmsta_10_i_0, C
         => \fsmsta[21]_net_1\, D => \fsmsta_nxt_9_m[21]\, Y => 
        \fsmsta_8[21]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_0\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_3_601_0_1, D => N_1717, Y => fsmsta_8_3_601_0);
    
    \framesync[2]\ : SLE
      port map(D => \framesync_7[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[2]_net_1\);
    
    \fsmmod_ns_0_a4[5]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => \pedetect\, B => \SCLSCL\, C => un115_fsmdet, 
        D => \fsmmod[1]_net_1\, Y => N_1058);
    
    \fsmmod_ns_0_a4[0]\ : CFG4
      generic map(INIT => x"AAA2")

      port map(A => \fsmmod[6]_net_1\, B => \starto_en\, C => 
        N_1040, D => N_64, Y => N_1048);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sersta_RNO[4]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => N_127, B => N_23, C => \sersta_32_i_a2_9[4]\, 
        D => \sersta_32_i_a2_7[4]\, Y => N_100_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_2_647_i_0_m2_0\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \COREI2C_0_2_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_120);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307_a3_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \ack\, B => N_2177, C => N_133, D => 
        fsmsta_8_28_307_a3_0_1, Y => N_1486);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_10[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[22]_net_1\, B => \fsmsta[21]_net_1\, 
        C => \COREI2C_0_2_INT[0]\, D => \sersta_32_i_a2_7[3]\, Y
         => \sersta_32_i_a2_10[3]\);
    
    un1_fsmsta_1_i_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => \fsmsta[15]_net_1\, B => \fsmsta[16]_net_1\, 
        Y => \un1_fsmsta_1_i_0_o2_0\);
    
    SDAO_int_1_sqmuxa_7 : CFG3
      generic map(INIT => x"47")

      port map(A => \nedetect\, B => un33_fsmsta, C => N_2177, Y
         => \SDAO_int_1_sqmuxa_7\);
    
    PCLK_count1_1_sqmuxa : CFG4
      generic map(INIT => x"00D0")

      port map(A => \PCLK_count1_ov_1_sqmuxa_1\, B => bclke, C
         => PCLK_count2_ov_6_1, D => \un1_PCLK_count1_0_sqmuxa\, 
        Y => \PCLK_count1_1_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_a6_0_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \framesync[3]_net_1\, B => 
        \framesync[0]_net_1\, Y => N_1658_1);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_5[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[1]_net_1\, Y
         => \sersta_32_i_a2_5[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3_0_1\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \ack\, B => \fsmsta[23]_net_1\, C => 
        \adrcompen\, D => \adrcomp\, Y => fsmsta_8_5_555_a3_0_1);
    
    \fsmsta[28]\ : SLE
      port map(D => \fsmsta_8[28]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[28]_net_1\);
    
    \serCON_WRITE_PROC.un16_fsmmod_0_a2_0_a3\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \sercon[4]_net_1\, B => \fsmmod[1]_net_1\, C
         => \fsmmod[6]_net_1\, Y => un16_fsmmod);
    
    \fsmsta_RNO_0[14]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \COREI2C_0_2_SDAO[0]\, B => N_2196, C => 
        N_2186, Y => N_36_i_1);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[2]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        PCLK_count2_ov_6_1, C => CO1, D => \PCLK_count1_1_sqmuxa\, 
        Y => \PCLK_count1_10[2]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns[16]\ : CFG4
      generic map(INIT => x"F808")

      port map(A => N_2177, B => \fsmsta[16]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_ns_1[16]\, Y => 
        \fsmsta_8[16]\);
    
    framesync_0_sqmuxa : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[6]_net_1\, C
         => un70_fsmsta, D => un19_framesync_1, Y => 
        \framesync_0_sqmuxa\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[2]\ : CFG3
      generic map(INIT => x"48")

      port map(A => CO1_0, B => PCLK_count2_ov_6_1, C => 
        \PCLK_count2[2]_net_1\, Y => \PCLK_count2_3[2]\);
    
    \sersta[1]\ : SLE
      port map(D => \sersta_32[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[1]_net_1\);
    
    \fsmdet[4]\ : SLE
      port map(D => N_859_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[4]_net_1\);
    
    \serDAT_WRITE_PROC.ack_7_u\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \SDAInt\, B => \ack\, C => 
        un1_serdat_2_sqmuxa_1_1, D => \serdat_0_sqmuxa\, Y => 
        ack_7);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_3\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[13]_net_1\, 
        C => \fsmsta[11]_net_1\, D => \fsmsta[10]_net_1\, Y => 
        un135_ens1_3);
    
    \fsmsync[7]\ : SLE
      port map(D => \fsmsync_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[7]_net_1\);
    
    \indelay[0]\ : SLE
      port map(D => N_57_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[0]_net_1\);
    
    \fsmsta[29]\ : SLE
      port map(D => \fsmsta_8[29]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[29]_net_1\);
    
    \fsmdet[0]\ : SLE
      port map(D => N_867_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[0]_net_1\);
    
    \fsmsta_RNO[13]\ : CFG4
      generic map(INIT => x"0D00")

      port map(A => N_2186, B => N_2177, C => un136_framesync, D
         => N_82, Y => N_34_i_0);
    
    \sercon[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[7]_net_1\);
    
    ack_bit : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => \ack_bit_1_sqmuxa\, ALn => MSS_READY, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ack_bit\);
    
    \fsmsta[2]\ : SLE
      port map(D => N_1604_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[2]_net_1\);
    
    \fsmdet[2]\ : SLE
      port map(D => N_863_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[2]_net_1\);
    
    \fsmdet_RNO[2]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \fsmdet[3]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_863_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_m0[0]\ : CFG4
      generic map(INIT => x"00FE")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => un149_framesync, D => \framesync_0_sqmuxa\, Y => 
        \framesync_7_m0[3]\);
    
    \framesync[1]\ : SLE
      port map(D => \framesync_7[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[1]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32[1]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \sersta_32_5[1]\, B => N_72_mux, C => 
        \sersta_32_4[1]\, Y => \sersta_32[1]\);
    
    \serDAT_WRITE_PROC.serdat_9[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un105_ens1, B => \ack\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(0), Y => \serdat_9[0]\);
    
    \sercon[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[0]_net_1\);
    
    \fsmsync[1]\ : SLE
      port map(D => N_976_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[1]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[27]\ : CFG4
      generic map(INIT => x"3320")

      port map(A => \un1_fsmsta_6\, B => un136_framesync, C => 
        \fsmsta_nxt_9_m_0[27]\, D => fsmsta_nxt_1_sqmuxa_24_s4_1, 
        Y => \fsmsta_8[27]\);
    
    \serDAT_WRITE_PROC.serdat_9[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(4), B => 
        un105_ens1, C => \serdat[3]_net_1\, Y => \serdat_9[4]\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_1_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        un57_fsmsta_1_0);
    
    \fsmmod[0]\ : SLE
      port map(D => N_1032_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[0]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_0_2[3]\ : CFG3
      generic map(INIT => x"28")

      port map(A => N_2179, B => \framesync[3]_net_1\, C => 
        N_1652, Y => N_161_2);
    
    SCLO_int_RNI9K79 : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_2_SCLO[0]\, Y => 
        COREI2C_0_2_SCLO_i(0));
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555\ : CFG4
      generic map(INIT => x"F0F4")

      port map(A => N_2177, B => fsmsta_8_5_555_a3_0_1, C => 
        N_1680, D => N_2181, Y => fsmsta_8_5_555_0);
    
    \fsmmod[6]\ : SLE
      port map(D => \fsmmod_ns[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[6]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_9[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \fsmsta[14]_net_1\, B => \fsmsta[6]_net_1\, C
         => \COREI2C_0_2_INT[0]\, D => \sersta_32_i_a2_6[4]\, Y
         => \sersta_32_i_a2_9[4]\);
    
    \sercon[4]\ : SLE
      port map(D => \sercon_9[4]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sercon[4]_net_1\);
    
    \FSMSYNC_SYNC_PROC.un139_ens1_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREI2C_0_2_INT[0]\, B => \SCLInt\, Y => 
        un139_ens1_0);
    
    adrcomp_2_sqmuxa_i_o2_0 : CFG4
      generic map(INIT => x"3F20")

      port map(A => seradr0apb(0), B => \ack\, C => 
        un13_adrcompen, D => \adrcomp_2_sqmuxa_i_a2_1_5\, Y => 
        N_2187);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_13_406\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \fsmsta[0]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1549);
    
    SCLO_int : SLE
      port map(D => un149_ens1_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_2_SCLO[0]\);
    
    \fsmmod[2]\ : SLE
      port map(D => N_1029_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[2]_net_1\);
    
    \sersta[3]\ : SLE
      port map(D => N_99_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sersta[3]_net_1\);
    
    \FRAMESYNC_WRITE_PROC.framesync_7[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \framesync_7_m0[3]\, B => framesync_7_sm0, Y
         => \framesync_7_m2[3]\);
    
    \serCON_WRITE_PROC.sercon_8_0_a3_1_0[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_2179, B => \sercon[6]_net_1\, Y => 
        \sercon_8_0_a3_1_0[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_28_307\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => \fsmsta[15]_net_1\, B => N_2177, C => N_2181, 
        D => N_1486, Y => N_1470);
    
    \fsmsync[6]\ : SLE
      port map(D => N_966_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[6]_net_1\);
    
    \SDAI_ff_reg[2]\ : SLE
      port map(D => \SDAI_ff_reg_4[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[2]_net_1\);
    
    \serdat_RNI9T7T[3]\ : CFG4
      generic map(INIT => x"03F5")

      port map(A => \COREI2C_0_2_INT[0]\, B => \serdat[3]_net_1\, 
        C => CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \PRDATA_3_1_1[3]\);
    
    \PCLK_count1[0]\ : SLE
      port map(D => \PCLK_count1_10[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[0]_net_1\);
    
    \fsmsta_RNO[17]\ : CFG4
      generic map(INIT => x"0B08")

      port map(A => \fsmsta[17]_net_1\, B => N_2177, C => N_2181, 
        D => N_2173_i_1, Y => N_2173_i_0);
    
    \fsmsync_ns_i_0_a2_0[2]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => \fsmsync[7]_net_1\, B => \fsmsync[6]_net_1\, 
        C => N_64, D => \fsmsync[5]_net_1\, Y => N_104);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_5_555_a3\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_2177, B => N_172, C => fsmsta_8_5_555_a3_0, 
        D => N_1622_2, Y => N_1680);
    
    \fsmsta_RNO[19]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_2199, B => un136_framesync, C => N_157, Y
         => N_2174_i_0);
    
    \fsmsync_ns_i_0_1_tz[3]\ : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \sercon[4]_net_1\, B => \fsmsync[5]_net_1\, C
         => N_130, D => un70_fsmsta, Y => 
        \fsmsync_ns_i_0_1_tz[3]_net_1\);
    
    \fsmsta[0]\ : SLE
      port map(D => N_1549, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[0]_net_1\);
    
    un1_fsmsta_6 : CFG3
      generic map(INIT => x"0E")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => N_2177, Y => \un1_fsmsta_6\);
    
    \serdat[3]\ : SLE
      port map(D => \serdat_9[3]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[3]_net_1\);
    
    \serCON_WRITE_PROC.un60_ens1_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \framesync[2]_net_1\, B => 
        \framesync[1]_net_1\, C => \framesync[0]_net_1\, Y => 
        N_1652);
    
    \fsmmod_ns_i_a4_1[2]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \COREI2C_0_2_INT[0]\, B => \sercon[5]_net_1\, 
        C => N_1041, D => \fsmmod_ns_i_a4_1_0[2]_net_1\, Y => 
        N_1054);
    
    \sersta_RNIM6MR1[2]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[5]\, C => \sersta[2]_net_1\, D => 
        \sercon[5]_net_1\, Y => N_1219);
    
    \serDAT_WRITE_PROC.serdat_9[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => 
        un105_ens1, C => \serdat[5]_net_1\, Y => \serdat_9[6]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_i_0\ : CFG4
      generic map(INIT => x"CFEE")

      port map(A => N_2182, B => N_2181, C => \fsmsta[9]_net_1\, 
        D => N_2177, Y => fsmsta_8_4_577_i_0);
    
    \fsmsta[5]\ : SLE
      port map(D => N_42_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[5]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2[0]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \COREI2C_0_2_INT[0]\, B => \fsmsta[9]_net_1\, 
        Y => \sersta_32_2[0]\);
    
    nedetect : SLE
      port map(D => \nedetect_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => rtn_i_0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \nedetect\);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => m7_3, B => fsmsta_8_20_379_i_0_a3_3, C => 
        \fsmsta[1]_net_1\, D => \fsmsta[11]_net_1\, Y => N_72_mux);
    
    adrcompen_2_sqmuxa_i : CFG4
      generic map(INIT => x"FFBA")

      port map(A => un16_fsmmod, B => N_2177, C => \nedetect\, D
         => \fsmdet[3]_net_1\, Y => adrcompen_2_sqmuxa_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_3[0]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \PCLK_count2[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, Y => 
        \PCLK_count2_3[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_1_676_i_0_m2\ : CFG3
      generic map(INIT => x"D1")

      port map(A => \COREI2C_0_2_SDAO[0]\, B => N_2177, C => 
        \fsmsta[12]_net_1\, Y => N_124);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl[1]\ : CFG4
      generic map(INIT => x"7B48")

      port map(A => CO0, B => framesync_7_e2, C => 
        \framesync[1]_net_1\, D => \fsmdet[3]_net_1\, Y => 
        \framesync_7[1]\);
    
    \serCON_WRITE_PROC.sercon_9[4]\ : CFG4
      generic map(INIT => x"F202")

      port map(A => \sercon_8_2[4]\, B => \fsmsta_cnst[0]\, C => 
        un5_penable, D => CoreAPB3_0_APBmslave0_PWDATA(4), Y => 
        \sercon_9[4]\);
    
    \fsmsta_RNO[14]\ : CFG4
      generic map(INIT => x"00B8")

      port map(A => \fsmsta[14]_net_1\, B => N_2177, C => 
        N_36_i_1, D => un136_framesync, Y => N_36_i_0);
    
    adrcomp_2_sqmuxa_i_o2_1_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[11]_net_1\, B => \fsmsta[10]_net_1\, 
        C => \fsmsta[6]_net_1\, D => \fsmsta[5]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_o2_1_3\);
    
    \indelay_RNO[1]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => \indelay[1]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_76, Y => N_55_i_0);
    
    \FSMSTA_SYNC_PROC.un133_framesync\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \pedetect\, B => \fsmsta[23]_net_1\, C => 
        un1_fsmmod, D => N_2177, Y => un133_framesync);
    
    \FSMSTA_SYNC_PROC.un136_framesync_0_o3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un133_framesync, B => N_2181, Y => 
        un136_framesync);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[0]\ : CFG4
      generic map(INIT => x"0048")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        PCLK_count2_ov_6_1, C => \un1_PCLK_count1_0_sqmuxa\, D
         => \PCLK_count1_1_sqmuxa\, Y => \PCLK_count1_10[0]\);
    
    \serDAT_WRITE_PROC.un92_fsmsta\ : CFG2
      generic map(INIT => x"2")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, Y => 
        un92_fsmsta);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[22]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \SDAInt\, B => \un1_fsmsta_6\, C => \ack\, Y
         => \fsmsta_nxt_9_m[22]\);
    
    \serDAT_WRITE_PROC.un134_fsmsta\ : CFG3
      generic map(INIT => x"10")

      port map(A => un57_fsmsta, B => \fsmdet[3]_net_1\, C => 
        un25_fsmsta, Y => un134_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_i_RNO\ : CFG4
      generic map(INIT => x"C010")

      port map(A => \nedetect\, B => \COREI2C_0_2_INT[0]\, C => 
        bsd7_i_m_0, D => un105_ens1, Y => bsd7_i_m);
    
    PCLK_count1_0_sqmuxa_1_1 : CFG4
      generic map(INIT => x"0111")

      port map(A => \sercon[0]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => 
        \PCLK_count1_0_sqmuxa_1_1\);
    
    \FRAMESYNC_WRITE_PROC.un19_framesync_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[13]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, Y => un19_framesync_1);
    
    adrcompen_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => un16_fsmmod, B => \fsmdet[3]_net_1\, Y => 
        \adrcompen_0_sqmuxa\);
    
    \serCON_WRITE_PROC.un70_ens1_i_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => mst, B => \adrcomp\, Y => N_2179);
    
    \fsmsync_ns_i_0_o2[3]\ : CFG3
      generic map(INIT => x"37")

      port map(A => N_67, B => \fsmsync[4]_net_1\, C => N_66, Y
         => N_63);
    
    \fsmsta[1]\ : SLE
      port map(D => N_1586_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[1]_net_1\);
    
    \fsmmod_ns_0_a4[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \nedetect\, B => un115_fsmdet, C => 
        \fsmmod[5]_net_1\, Y => N_1050);
    
    \framesync[0]\ : SLE
      port map(D => \framesync_7[0]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \framesync[0]_net_1\);
    
    \un2_framesync_1_1.CO0\ : CFG3
      generic map(INIT => x"08")

      port map(A => \nedetect\, B => \framesync[0]_net_1\, C => 
        un70_fsmsta, Y => CO0);
    
    bsd7_tmp : SLE
      port map(D => bsd7_tmp_6, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7_tmp\);
    
    \fsmdet[3]\ : SLE
      port map(D => N_861_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[3]_net_1\);
    
    PCLKint_ff : SLE
      port map(D => PCLKint_ff_2, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint_ff\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_23_351_i_0_1\ : CFG4
      generic map(INIT => x"3AFF")

      port map(A => \COREI2C_0_2_SDAO[0]\, B => 
        \fsmsta[20]_net_1\, C => N_2177, D => N_2178, Y => 
        fsmsta_8_23_351_i_0_1);
    
    \serdat[6]\ : SLE
      port map(D => \serdat_9[6]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[6]_net_1\);
    
    \fsmmod_ns_i_o3_1[2]\ : CFG2
      generic map(INIT => x"7")

      port map(A => un70_fsmsta, B => \fsmmod[4]_net_1\, Y => 
        N_1041);
    
    \fsmmod_ns_0_o3_0_0[3]\ : CFG3
      generic map(INIT => x"B7")

      port map(A => \PCLKint\, B => \SCLInt\, C => \PCLKint_ff\, 
        Y => N_1034);
    
    \fsmdet_RNO[0]\ : CFG4
      generic map(INIT => x"E0A0")

      port map(A => \fsmdet[1]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SCLInt\, D => \SDAInt\, Y => N_867_i_0);
    
    \fsmmod_RNO[2]\ : CFG4
      generic map(INIT => x"0045")

      port map(A => N_1064, B => \fsmmod[2]_net_1\, C => N_1046, 
        D => un115_fsmdet, Y => N_1029_i_0);
    
    \serCON_WRITE_PROC.un5_penable\ : CFG3
      generic map(INIT => x"80")

      port map(A => un3_penable_1, B => un5_penable_1, C => N_40, 
        Y => un5_penable);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[5]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \fsmsta[5]_net_1\, B => \SDAInt\, C => N_2171, 
        Y => N_80);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[24]\ : CFG4
      generic map(INIT => x"0805")

      port map(A => N_2177, B => \fsmsta[24]_net_1\, C => 
        un136_framesync, D => \fsmsta_8_1[24]\, Y => 
        \fsmsta_8[24]\);
    
    un1_PCLK_count1_0_sqmuxa_1_0 : CFG4
      generic map(INIT => x"08AF")

      port map(A => CO2, B => bclke, C => \PCLK_count1[3]_net_1\, 
        D => \sercon[7]_net_1\, Y => 
        \un1_PCLK_count1_0_sqmuxa_1_0\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[16]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[16]\);
    
    starto_en_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \fsmmod[1]_net_1\, B => N_64, C => \busfree\, 
        D => \SCLInt\, Y => N_60);
    
    \fsmmod_ns_0_o3_0[3]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \sercon[4]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => \sercon[5]_net_1\, Y => N_1040);
    
    \serDAT_WRITE_PROC.serdat_9[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(3), B => 
        un105_ens1, C => \serdat[2]_net_1\, Y => \serdat_9[3]\);
    
    bsd7 : SLE
      port map(D => bsd7_9_iv_i_0, CLK => FAB_CCC_GL0, EN => 
        \sercon[6]_net_1\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \bsd7\);
    
    PCLKint : SLE
      port map(D => PCLKint_3, CLK => FAB_CCC_GL0, EN => 
        un1_pclkint4_i_0, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLKint\);
    
    \PCLK_count1[1]\ : SLE
      port map(D => \PCLK_count1_10[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[1]_net_1\);
    
    \fsmsta[13]\ : SLE
      port map(D => N_34_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[13]_net_1\);
    
    \serdat[5]\ : SLE
      port map(D => \serdat_9[5]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[5]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1\ : CFG4
      generic map(INIT => x"4440")

      port map(A => un16_fsmmod, B => PCLK_count2_ov_6_0_a2_1_3, 
        C => \SCLInt\, D => PCLK_count2_ov_6_0_a2_1_4_tz, Y => 
        PCLK_count2_ov_6_1);
    
    \serDAT_WRITE_PROC.serdat_9[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        un105_ens1, C => \serdat[6]_net_1\, Y => \serdat_9[7]\);
    
    \sersta_RNIQAMR1[3]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[6]\, C => \sersta[3]_net_1\, D => 
        \sercon[6]_net_1\, Y => N_1220);
    
    \sersta_RNII2MR1[1]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[4]\, C => \sersta[1]_net_1\, D => 
        seradr0apb(4), Y => N_1218);
    
    un1_counter_rst_3 : CFG2
      generic map(INIT => x"B")

      port map(A => \PCLK_count1_1_sqmuxa\, B => 
        PCLK_count2_ov_6_1, Y => \un1_counter_rst_3\);
    
    \fsmsync_RNO[4]\ : CFG4
      generic map(INIT => x"0155")

      port map(A => N_1002, B => \fsmsync_ns_i_0_1_tz[3]_net_1\, 
        C => \COREI2C_0_2_INT[0]\, D => N_63, Y => N_970_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => N_2177);
    
    \SDAI_ff_reg[0]\ : SLE
      port map(D => \SDAI_ff_reg_4[0]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[0]_net_1\);
    
    \fsmsync_RNO[5]\ : CFG4
      generic map(INIT => x"0103")

      port map(A => \fsmsync[7]_net_1\, B => N_104, C => N_1002, 
        D => N_86, Y => N_968_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m2[13]\ : CFG4
      generic map(INIT => x"CACC")

      port map(A => \COREI2C_0_2_SDAO[0]\, B => 
        \fsmsta[13]_net_1\, C => N_2177, D => N_2196, Y => N_82);
    
    \fsmsta_RNO[12]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_1656, B => N_2186, C => N_2181, D => N_124, 
        Y => N_1774_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_o3_i_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \SDAInt\, B => \COREI2C_0_2_SDAO[0]\, Y => 
        N_172);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6_m1\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(7), B => 
        \serdat_0_sqmuxa\, Y => bsd7_tmp_6_m1);
    
    \serdat_RNIBV7T[4]\ : CFG4
      generic map(INIT => x"0F53")

      port map(A => \serdat[4]_net_1\, B => \sercon[4]_net_1\, C
         => CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[4]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => fsmsta_8_20_379_i_0_a3_3_0, B => 
        fsmsta_8_20_379_i_0_a3_3, C => N_2177, D => 
        fsmsta_8_20_379_i_0_a3_4, Y => N_145);
    
    adrcomp : SLE
      port map(D => N_2176_i_0, CLK => FAB_CCC_GL0, EN => 
        adrcomp_2_sqmuxa_i_0_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcomp\);
    
    \fsmsync_ns_0_0[0]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => N_70, B => \fsmsync_ns_0_0_1[0]_net_1\, C => 
        \fsmsync[7]_net_1\, D => \SCLInt\, Y => \fsmsync_ns[0]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601_m4\ : CFG4
      generic map(INIT => x"3074")

      port map(A => \fsmmod[0]_net_1\, B => \fsmdet[3]_net_1\, C
         => \fsmdet[1]_net_1\, D => \fsmmod[5]_net_1\, Y => 
        N_1717);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_5\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[18]_net_1\, B => \fsmsta[17]_net_1\, 
        C => un135_ens1_2, Y => un135_ens1_5);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[23]_net_1\, B => \fsmsta[7]_net_1\, Y
         => fsmsta_8_20_379_i_0_a3_3);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[11]_net_1\, 
        C => \fsmsta[10]_net_1\, D => \fsmsta[9]_net_1\, Y => 
        \sersta_32_i_a2_7[4]\);
    
    \SDAO_INT_WRITE_PROC.un25_fsmsta_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[15]_net_1\, 
        C => \fsmsta[18]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        un25_fsmsta_2);
    
    \sersta_RNIEULR1[0]\ : CFG4
      generic map(INIT => x"B391")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \PRDATA_3_1_1[3]\, C => \sersta[0]_net_1\, D => 
        seradr0apb(3), Y => N_1217);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_4_577_a3_0_2_0_i_o3_0\ : CFG4
      generic map(INIT => x"F4F0")

      port map(A => \PCLKint\, B => \PCLKint_ff\, C => N_1586_1, 
        D => \fsmmod[2]_net_1\, Y => N_2181);
    
    \fsmsta[17]\ : SLE
      port map(D => N_2173_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[17]_net_1\);
    
    \fsmmod_ns_i_o3[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_1041, B => N_997, Y => N_1046);
    
    adrcompen : SLE
      port map(D => \adrcompen_0_sqmuxa\, CLK => FAB_CCC_GL0, EN
         => adrcompen_2_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \adrcompen\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[26]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[26]\);
    
    \indelay[3]\ : SLE
      port map(D => N_51_i_0, CLK => FAB_CCC_GL0, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \indelay[3]_net_1\);
    
    \SDAI_ff_reg[1]\ : SLE
      port map(D => \SDAI_ff_reg_4[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SDAI_ff_reg[1]_net_1\);
    
    \fsmsta[8]\ : SLE
      port map(D => fsmsta_8_5_555_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[8]_net_1\);
    
    \fsmsync_ns_i_0_a2[5]\ : CFG3
      generic map(INIT => x"0D")

      port map(A => \fsmsync[5]_net_1\, B => N_64, C => 
        \fsmsync[2]_net_1\, Y => N_130);
    
    \ADRCOMP_WRITE_PROC.un20_adrcompen_i_0_o3\ : CFG2
      generic map(INIT => x"7")

      port map(A => un13_adrcompen, B => seradr0apb(0), Y => 
        N_133);
    
    \fsmdet[6]\ : SLE
      port map(D => SCLInt_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[6]_net_1\);
    
    \fsmsta_RNO[6]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \fsmsta[6]_net_1\, B => \SDAInt\, C => N_2171, 
        D => un136_framesync, Y => N_44_i_0);
    
    \fsmmod_ns_0[1]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1050, Y => \fsmmod_ns[1]\);
    
    ack_bit_1_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \COREI2C_0_2_INT[0]\, B => \sercon[6]_net_1\, 
        C => un134_fsmsta, D => un5_penable, Y => 
        \ack_bit_1_sqmuxa\);
    
    \fsmsync_ns_i_0_o2_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_70, B => \SCLInt\, Y => N_86);
    
    \FSMSTA_SYNC_PROC.un133_framesync_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \adrcomp\, B => \adrcompen\, Y => un1_fsmmod);
    
    pedetect_0_sqmuxa : CFG4
      generic map(INIT => x"2000")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \pedetect_0_sqmuxa\);
    
    mst_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmmod[1]_net_1\, B => \fsmmod[6]_net_1\, Y
         => mst);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[28]_net_1\, B => \fsmsta[29]_net_1\, 
        C => un57_fsmsta_1_0, D => un57_fsmsta_0, Y => 
        un57_fsmsta);
    
    \fsmsta_RNO[11]\ : CFG3
      generic map(INIT => x"10")

      port map(A => N_2181, B => fsmsta_8_2_647_i_0_0, C => 
        N_1656, Y => N_1751_i_0);
    
    \PRDATA_1[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \sercon[1]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => \serdat[1]_net_1\, Y
         => N_1197);
    
    PCLK_count1_0_sqmuxa_3 : CFG4
      generic map(INIT => x"4CCC")

      port map(A => \PCLK_count1[1]_net_1\, B => 
        \un1_pclk_count191\, C => \PCLK_count1[3]_net_1\, D => 
        \PCLK_count1[2]_net_1\, Y => \PCLK_count1_0_sqmuxa_3\);
    
    adrcomp_2_sqmuxa_i_a3_4 : CFG4
      generic map(INIT => x"0800")

      port map(A => \sercon[2]_net_1\, B => \adrcompen\, C => 
        \framesync[3]_net_1\, D => \adrcomp_2_sqmuxa_i_a3_3\, Y
         => \adrcomp_2_sqmuxa_i_a3_4\);
    
    \serSTA_WRITE_PROC.sersta_32_4[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[16]_net_1\, B => \fsmsta[8]_net_1\, C
         => \fsmsta[20]_net_1\, D => \fsmsta[2]_net_1\, Y => 
        \sersta_32_4[1]\);
    
    SDAO_int_RNIV27C : CFG1
      generic map(INIT => "01")

      port map(A => \COREI2C_0_2_SDAO[0]\, Y => 
        COREI2C_0_2_SDAO_i(0));
    
    un1_PCLK_count1_0_sqmuxa : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \PCLK_count1_0_sqmuxa_4\, B => 
        \PCLK_count1_0_sqmuxa_3\, C => 
        \un1_PCLK_count1_0_sqmuxa_0\, D => 
        \un1_PCLK_count1_0_sqmuxa_1_0\, Y => 
        \un1_PCLK_count1_0_sqmuxa\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8[22]\ : CFG4
      generic map(INIT => x"3222")

      port map(A => \fsmsta_nxt_9_m[22]\, B => un136_framesync, C
         => \fsmsta[22]_net_1\, D => N_2177, Y => \fsmsta_8[22]\);
    
    \sersta[4]\ : SLE
      port map(D => N_100_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[4]_net_1\);
    
    SCLInt : SLE
      port map(D => \SCLI_ff_reg[0]_net_1\, CLK => FAB_CCC_GL0, 
        EN => un1_rtn_3_1, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \SCLInt\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[1]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[0]_net_1\, B => 
        \PCLK_count1[1]_net_1\, C => \un1_counter_rst_3\, D => 
        \un1_PCLK_count1_0_sqmuxa\, Y => \PCLK_count1_10[1]\);
    
    \serdat_RNI6TF21[7]\ : CFG4
      generic map(INIT => x"503F")

      port map(A => seradr0apb(7), B => \serdat[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => \PRDATA_3_1_1[7]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1_4\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[6]_net_1\, B => \fsmsta[12]_net_1\, C
         => \fsmsta[9]_net_1\, D => \fsmsta[5]_net_1\, Y => 
        un135_ens1_4);
    
    \fsmsync_ns_0_0_o2[0]\ : CFG3
      generic map(INIT => x"F4")

      port map(A => \fsmmod[1]_net_1\, B => N_117_1, C => N_64, Y
         => N_70);
    
    \fsmmod_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \nedetect\, B => \fsmmod[3]_net_1\, C => 
        un115_fsmdet, D => N_1060, Y => N_1032_i_0);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \bsd7_tmp\, B => \SCLInt\, C => 
        \COREI2C_0_2_INT[0]\, D => un57_fsmsta, Y => 
        bsd7_tmp_i_m_2);
    
    \fsmsta[11]\ : SLE
      port map(D => N_1751_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[11]_net_1\);
    
    un1_serdat_2_sqmuxa : CFG4
      generic map(INIT => x"F0F8")

      port map(A => \sercon[6]_net_1\, B => \pedetect\, C => 
        un105_ens1, D => \un1_serdat_2_sqmuxa_1_0\, Y => 
        \un1_serdat_2_sqmuxa_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_RNIEH881\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \nedetect\, B => \COREI2C_0_2_INT[0]\, C => 
        un57_fsmsta, D => un105_ens1, Y => bsd7_tmp_6_sn_N_10_mux);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[1]_net_1\, Y => \SDAI_ff_reg_4[2]\);
    
    \INDELAY_WRITE_PROC.indelay_4_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \indelay[1]_net_1\, B => \indelay[3]_net_1\, 
        Y => N_66);
    
    PCLK_count2_ov : SLE
      port map(D => PCLK_count2_ov_6, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2_ov\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_0[25]\ : CFG4
      generic map(INIT => x"55CF")

      port map(A => \fsmsta[25]_net_1\, B => \SDAInt\, C => 
        un57_fsmsta_1_0, D => N_2177, Y => \fsmsta_8_i_0[25]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO[27]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \SDAInt\, B => \ack\, Y => 
        \fsmsta_nxt_9_m_0[27]\);
    
    \fsmsta[26]\ : SLE
      port map(D => \fsmsta_8[26]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[26]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_2_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[5]_net_1\, B => \fsmsta[13]_net_1\, Y
         => N_127);
    
    \fsmsync_RNO[2]\ : CFG3
      generic map(INIT => x"04")

      port map(A => N_1002, B => \COREI2C_0_2_INT[0]\, C => N_130, 
        Y => N_974_i_0);
    
    \sercon[3]\ : SLE
      port map(D => \sercon_9[3]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREI2C_0_2_INT[0]\);
    
    \fsmsync_ns_i_0_o2_0[4]\ : CFG4
      generic map(INIT => x"FF7F")

      port map(A => \indelay[2]_net_1\, B => \indelay[0]_net_1\, 
        C => \fsmsync[4]_net_1\, D => N_66, Y => N_84);
    
    \BUSFREE_WRITE_PROC.un105_fsmdet\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \sercon[6]_net_1\, B => N_1586_1, C => 
        un16_fsmmod, D => N_1064, Y => un105_fsmdet);
    
    \fsmmod[5]\ : SLE
      port map(D => \fsmmod_ns[1]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[5]_net_1\);
    
    un1_serdat_2_sqmuxa_1 : CFG4
      generic map(INIT => x"0C08")

      port map(A => un92_fsmsta, B => \pedetect\, C => un105_ens1, 
        D => \un1_serdat40\, Y => un1_serdat_2_sqmuxa_1_1);
    
    \fsmdet[5]\ : SLE
      port map(D => N_857_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmdet[5]_net_1\);
    
    \fsmmod[1]\ : SLE
      port map(D => \fsmmod_ns[5]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmmod[1]_net_1\);
    
    \fsmdet_RNO[4]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[6]_net_1\, B => \fsmdet[4]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_859_i_0);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_o4_0\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => \framesync[3]_net_1\, B => \bsd7\, C => 
        un57_fsmsta, D => un70_fsmsta, Y => N_1465);
    
    \fsmdet_RNO[1]\ : CFG4
      generic map(INIT => x"E000")

      port map(A => \fsmdet[4]_net_1\, B => \fsmdet[2]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_865_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_3_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[27]_net_1\, B => \fsmsta[26]_net_1\, 
        C => \fsmsta[25]_net_1\, D => \fsmsta[24]_net_1\, Y => 
        fsmsta_8_20_379_i_0_a3_3_0);
    
    \serSTA_WRITE_PROC.sersta_32_4[2]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsta[9]_net_1\, B => \fsmsta[23]_net_1\, C
         => \fsmsta[10]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_4[2]\);
    
    \fsmsync[4]\ : SLE
      port map(D => N_970_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[4]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_3_601\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[10]_net_1\, C => 
        N_1657_2, D => fsmsta_8_3_601_0, Y => N_1701);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a2_0\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_172, B => N_2182, C => N_2193, Y => N_165);
    
    \fsmsta[14]\ : SLE
      port map(D => N_36_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[14]_net_1\);
    
    \fsmsync_ns_i_a3_1_0_a2[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmmod[4]_net_1\, B => \fsmmod[5]_net_1\, C
         => \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\, Y => N_1002);
    
    SCLSCL_1_sqmuxa_i : CFG2
      generic map(INIT => x"D")

      port map(A => \fsmmod[1]_net_1\, B => \pedetect\, Y => 
        SCLSCL_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[27]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[27]_net_1\, C => N_172, 
        Y => fsmsta_nxt_1_sqmuxa_24_s4_1);
    
    \fsmsta_RNO[3]\ : CFG4
      generic map(INIT => x"00BF")

      port map(A => \framesync[0]_net_1\, B => 
        fsmsta_8_10_476_i_a6_0, C => N_1624, D => 
        fsmsta_8_10_476_i_1, Y => N_1622_i_0);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \serdat[6]_net_1\, B => \serdat[5]_net_1\, C
         => \serdat[4]_net_1\, D => \serdat[3]_net_1\, Y => 
        un13_adrcompen_4);
    
    \sercon[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[5]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un57_fsmsta_0\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \fsmsta[7]_net_1\, B => \fsmsta[9]_net_1\, C
         => \fsmsta[8]_net_1\, Y => un57_fsmsta_0);
    
    \PRDATA_3[2]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        seradr0apb(2), C => N_1198, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_1216);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_RNO_0[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_2177, B => \fsmsta[26]_net_1\, C => N_172, 
        Y => fsmsta_nxt_1_sqmuxa_18_s5_1);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_enl_ns_1[3]\ : CFG4
      generic map(INIT => x"7F80")

      port map(A => \framesync[1]_net_1\, B => 
        \framesync[2]_net_1\, C => CO0, D => \framesync[3]_net_1\, 
        Y => \framesync_7_enl_ns_1[3]\);
    
    \serDAT_WRITE_PROC.serdat_9[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        un105_ens1, C => \serdat[4]_net_1\, Y => \serdat_9[5]\);
    
    nedetect_RNO : CFG3
      generic map(INIT => x"7F")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_i_0);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_4_tz\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[1]_net_1\, C
         => \COREI2C_0_2_SCLO[0]\, D => \busfree\, Y => 
        PCLK_count2_ov_6_0_a2_1_4_tz);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_10_476_i_o6_0\ : CFG4
      generic map(INIT => x"3430")

      port map(A => \fsmsta[23]_net_1\, B => \framesync[3]_net_1\, 
        C => N_1586_1, D => un1_fsmmod, Y => N_1624);
    
    serdat_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => un92_fsmsta, B => \COREI2C_0_2_INT[0]\, Y => 
        \serdat_0_sqmuxa\);
    
    \fsmsta[9]\ : SLE
      port map(D => N_2172_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[9]_net_1\);
    
    \SDAO_INT_WRITE_PROC.un70_fsmsta\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \framesync[0]_net_1\, B => 
        \framesync[3]_net_1\, C => \framesync[2]_net_1\, D => 
        \framesync[1]_net_1\, Y => un70_fsmsta);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1_RNO\ : CFG3
      generic map(INIT => x"02")

      port map(A => un57_fsmsta, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => 
        \COREI2C_0_2_INT[0]\, Y => \PWDATA_i_m_1[7]\);
    
    \fsmsta[25]\ : SLE
      port map(D => N_2175_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[25]_net_1\);
    
    \fsmmod_RNO[4]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => N_1046, B => N_1054, C => 
        \fsmmod_ns_i_0[2]_net_1\, D => un115_fsmdet, Y => 
        N_1026_i_0);
    
    \fsmsta[12]\ : SLE
      port map(D => N_1774_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[12]_net_1\);
    
    \CLK_COUNTER1_PROC.un12_pclk_count1_1.CO3\ : CFG4
      generic map(INIT => x"777F")

      port map(A => \PCLK_count1[3]_net_1\, B => 
        \PCLK_count1[2]_net_1\, C => \PCLK_count1[1]_net_1\, D
         => \PCLK_count1[0]_net_1\, Y => un12_pclk_count1);
    
    adrcomp_RNO : CFG3
      generic map(INIT => x"15")

      port map(A => \adrcomp_2_sqmuxa_i_0_0_0\, B => 
        \COREI2C_0_2_INT[0]\, C => N_2192, Y => N_2176_i_0);
    
    \SCLI_ff_reg[2]\ : SLE
      port map(D => \SCLI_ff_reg_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SCLI_ff_reg[2]_net_1\);
    
    \fsmsync_RNO[3]\ : CFG4
      generic map(INIT => x"0405")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => N_972_i_0);
    
    \fsmsync[3]\ : SLE
      port map(D => N_972_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[3]_net_1\);
    
    \serCON_WRITE_PROC.sercon_8_0_1[3]\ : CFG4
      generic map(INIT => x"AAEA")

      port map(A => N_163, B => \sercon_8_0_a3_1_0[3]\, C => 
        \pedetect\, D => N_2177, Y => \sercon_8_0_1[3]\);
    
    \PCLK_count2[1]\ : SLE
      port map(D => \PCLK_count2_3[1]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[1]_net_1\);
    
    PCLKint_ff_RNIFJ191 : CFG3
      generic map(INIT => x"20")

      port map(A => \fsmmod[2]_net_1\, B => \PCLKint\, C => 
        \PCLKint_ff\, Y => \fsmsta_cnst[0]\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2_1_3\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsync[2]_net_1\, B => \fsmdet[1]_net_1\, C
         => \fsmdet[3]_net_1\, D => PCLK_count2_ov_6_0_a2_1_0, Y
         => PCLK_count2_ov_6_0_a2_1_3);
    
    \fsmsta[20]\ : SLE
      port map(D => N_1520_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[20]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_7[2]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[26]_net_1\, B => \fsmsta[18]_net_1\, 
        C => \COREI2C_0_2_INT[0]\, D => \sersta_32_4[2]\, Y => 
        \sersta_32_7[2]\);
    
    busfree : SLE
      port map(D => \fsmdet_i_0[3]\, CLK => FAB_CCC_GL0, EN => 
        un105_fsmdet, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \busfree\);
    
    \PCLK_count1[2]\ : SLE
      port map(D => \PCLK_count1_10[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count1[2]_net_1\);
    
    \fsmmod_ns_0_a4_0_4_2[3]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \fsmsta[29]_net_1\, B => \PCLKint_ff\, C => 
        \PCLKint\, D => \fsmsta[28]_net_1\, Y => 
        \fsmmod_ns_0_a4_0_4_2[3]_net_1\);
    
    \fsmsync_ns_i_1[6]\ : CFG4
      generic map(INIT => x"F7F4")

      port map(A => \SDAInt\, B => \fsmsync[1]_net_1\, C => 
        N_1002, D => N_997, Y => \fsmsync_ns_i_1[6]_net_1\);
    
    adrcomp_2_sqmuxa_i_a2_1_2 : CFG4
      generic map(INIT => x"8421")

      port map(A => seradr0apb(6), B => seradr0apb(5), C => 
        \serdat[5]_net_1\, D => \serdat[4]_net_1\, Y => 
        \adrcomp_2_sqmuxa_i_a2_1_2\);
    
    \sercon[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un5_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sercon[6]_net_1\);
    
    SDAO_int : SLE
      port map(D => N_1449, CLK => FAB_CCC_GL0, EN => 
        SDAO_int_1_sqmuxa_i_0, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \COREI2C_0_2_SDAO[0]\);
    
    \fsmsta[18]\ : SLE
      port map(D => \fsmsta_8[18]\, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[18]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[19]_net_1\, B => \fsmsta[20]_net_1\, 
        C => \fsmsta[16]_net_1\, D => \fsmsta[18]_net_1\, Y => 
        \sersta_32_i_a2_7[3]\);
    
    \fsmsta_RNO[23]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => N_145, B => N_2181, C => N_166, D => 
        fsmsta_8_20_379_i_0_o2_0, Y => N_1543_i_0);
    
    \FRAMESYNC_WRITE_PROC.framesync_7_e2\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \nedetect\, B => un70_fsmsta, C => N_2177, D
         => framesync_7_sm0, Y => framesync_7_e2);
    
    \fsmsync_ns_0_0_1[0]\ : CFG4
      generic map(INIT => x"F8FA")

      port map(A => \SCLInt\, B => \fsmsync[3]_net_1\, C => 
        N_1002, D => N_84, Y => \fsmsync_ns_0_0_1[0]_net_1\);
    
    \serSTA_WRITE_PROC.sersta_32_i_a2_8[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta[15]_net_1\, C
         => \fsmsta[6]_net_1\, D => \fsmsta[17]_net_1\, Y => 
        \sersta_32_i_a2_8[3]\);
    
    \ADRCOMP_WRITE_PROC.un13_adrcompen\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \serdat[2]_net_1\, B => \serdat[1]_net_1\, C
         => \serdat[0]_net_1\, D => un13_adrcompen_4, Y => 
        un13_adrcompen);
    
    \serSTA_WRITE_PROC.sersta_31_4_0_.m22\ : CFG2
      generic map(INIT => x"1")

      port map(A => \fsmsta[4]_net_1\, B => \fsmsta[0]_net_1\, Y
         => N_23);
    
    \SDAINT_WRITE_PROC.SDAI_ff_reg_4[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sercon[6]_net_1\, B => 
        \SDAI_ff_reg[0]_net_1\, Y => \SDAI_ff_reg_4[1]\);
    
    \fsmsta_RNO[2]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \fsmsta[2]_net_1\, B => \fsmsta_cnst[0]\, C
         => N_1586_1, D => N_1656, Y => N_1604_i_0);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1_RNINIE91 : CFG4
      generic map(INIT => x"FC54")

      port map(A => \un1_ens1_pre_1_sqmuxa_0_a2_1\, B => 
        \pedetect\, C => un136_framesync, D => N_161_2, Y => 
        un1_ens1_pre_1_sqmuxa_i_0);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \fsmsta_cnst[0]\, B => \adrcomp\, C => 
        fsmsta_8_9_509_0_1, D => N_1717, Y => fsmsta_8_9_509_0);
    
    \fsmsta_RNO[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => N_126, B => N_80, C => un136_framesync, Y => 
        N_42_i_0);
    
    \fsmsta[19]\ : SLE
      port map(D => N_2174_i_0, CLK => FAB_CCC_GL0, EN => 
        un1_ens1_pre_1_sqmuxa_i_0, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \fsmsta[19]_net_1\);
    
    \serDAT_WRITE_PROC.bsd7_9_iv_1\ : CFG4
      generic map(INIT => x"FBF8")

      port map(A => \PWDATA_i_m_1[7]\, B => un105_ens1, C => 
        \fsmdet[3]_net_1\, D => bsd7_tmp_i_m_2, Y => bsd7_9_iv_1);
    
    \fsmmod_ns_i_a4_1_0[2]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \fsmsta[29]_net_1\, B => \PCLKint_ff\, C => 
        \PCLKint\, D => \fsmsta[28]_net_1\, Y => 
        \fsmmod_ns_i_a4_1_0[2]_net_1\);
    
    \CLK_COUNT2_WRITE_PROC.PCLK_count2_ov_6_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \un1_pclk_count1_ov_1\, B => 
        PCLK_count2_ov_6_1, C => \PCLK_count1_ov\, D => 
        \un1_pclk_count1_ov\, Y => PCLK_count2_ov_6);
    
    \sersta_RNIUEMR1[4]\ : CFG4
      generic map(INIT => x"7632")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \PRDATA_3_1_1[7]\, C => \sersta[4]_net_1\, D => 
        \sercon[7]_net_1\, Y => N_1221);
    
    \fsmsync_ns_i_o3_0[6]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => un70_fsmsta, B => \fsmsync[5]_net_1\, C => 
        N_64, Y => N_995);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_20_379_i_0_a3_4\ : CFG3
      generic map(INIT => x"10")

      port map(A => \fsmsta[29]_net_1\, B => \fsmsta[28]_net_1\, 
        C => N_153_1, Y => fsmsta_8_20_379_i_0_a3_4);
    
    \PCLK_count2[2]\ : SLE
      port map(D => \PCLK_count2_3[2]\, CLK => FAB_CCC_GL0, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PCLK_count2[2]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_9_509\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1732, B => \fsmsta[4]_net_1\, C => N_1657_2, 
        D => fsmsta_8_9_509_0, Y => N_1631);
    
    \fsmmod_ns_0[3]\ : CFG4
      generic map(INIT => x"5444")

      port map(A => un115_fsmdet, B => 
        \fsmmod_ns_0_a4_0_4[3]_net_1\, C => \fsmmod[3]_net_1\, D
         => N_1034, Y => \fsmmod_ns[3]\);
    
    \fsmdet_RNO[6]\ : CFG1
      generic map(INIT => "01")

      port map(A => \SCLInt\, Y => SCLInt_i_0);
    
    \serSTA_WRITE_PROC.sersta_32[0]\ : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \sersta_32_2[0]\, B => N_72_mux, C => N_127, 
        D => \sersta_32_3[0]\, Y => \sersta_32[0]\);
    
    \FSMSYNC_SYNC_PROC.un135_ens1\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un135_ens1_4, B => \un1_fsmsta_1_i_0_o2_0\, C
         => un135_ens1_5, D => un135_ens1_3, Y => un135_ens1);
    
    un1_pclk_count1_ov_1_1 : CFG4
      generic map(INIT => x"1333")

      port map(A => \PCLK_count2[1]_net_1\, B => 
        \sercon[0]_net_1\, C => \PCLK_count2[3]_net_1\, D => 
        \PCLK_count2[2]_net_1\, Y => \un1_pclk_count1_ov_1_1\);
    
    \serdat[1]\ : SLE
      port map(D => \serdat_9[1]\, CLK => FAB_CCC_GL0, EN => 
        \un1_serdat_2_sqmuxa_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \serdat[1]_net_1\);
    
    SDAO_int_1_sqmuxa_3 : CFG4
      generic map(INIT => x"0301")

      port map(A => \fsmmod[6]_net_1\, B => \fsmmod[2]_net_1\, C
         => \fsmmod[0]_net_1\, D => \adrcomp\, Y => 
        \SDAO_int_1_sqmuxa_3\);
    
    \SDAO_INT_WRITE_PROC.SDAO_int_7_0_275_m5\ : CFG4
      generic map(INIT => x"7F40")

      port map(A => \ack_bit\, B => un33_fsmsta, C => un25_fsmsta, 
        D => N_1465, Y => N_1466);
    
    un1_serdat_2_sqmuxa_1_0 : CFG4
      generic map(INIT => x"00EF")

      port map(A => \fsmdet[3]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => un57_fsmsta, D => \un1_serdat40\, Y => 
        \un1_serdat_2_sqmuxa_1_0\);
    
    \serDAT_WRITE_PROC.bsd7_tmp_6\ : CFG4
      generic map(INIT => x"CFCA")

      port map(A => \bsd7_tmp\, B => bsd7_tmp_6_m1, C => 
        bsd7_tmp_6_sm0, D => bsd7_tmp_6_sn_N_10_mux, Y => 
        bsd7_tmp_6);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_a3[19]\ : CFG4
      generic map(INIT => x"0322")

      port map(A => un57_fsmsta_1_0, B => N_2177, C => \SDAInt\, 
        D => N_2178, Y => N_157);
    
    un1_pclk_count191 : CFG3
      generic map(INIT => x"4C")

      port map(A => \sercon[0]_net_1\, B => \sercon[7]_net_1\, C
         => \sercon[1]_net_1\, Y => \un1_pclk_count191\);
    
    \serDAT_WRITE_PROC.un105_ens1\ : CFG3
      generic map(INIT => x"80")

      port map(A => un3_penable_1, B => un105_ens1_1, C => N_40, 
        Y => un105_ens1);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, Y => \SCLI_ff_reg_3[2]\);
    
    \SCLINT_WRITE_PROC.SCLI_ff_reg_3[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => \sercon[6]_net_1\, B => 
        \SCLI_ff_reg[0]_net_1\, Y => \SCLI_ff_reg_3[1]\);
    
    \or_br.rtn_1\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => rtn_1);
    
    \fsmsync_ns_i_a3_1_0_a2_2[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \fsmmod[2]_net_1\, B => \fsmmod[3]_net_1\, C
         => \fsmmod[1]_net_1\, D => \fsmmod[0]_net_1\, Y => 
        \fsmsync_ns_i_a3_1_0_a2_2[2]_net_1\);
    
    un1_ens1_pre_1_sqmuxa_0_a2_1 : CFG4
      generic map(INIT => x"0D00")

      port map(A => un74_ens1, B => \COREI2C_0_2_INT[0]\, C => 
        N_1622_2, D => N_1586_1, Y => 
        \un1_ens1_pre_1_sqmuxa_0_a2_1\);
    
    \fsmdet_RNO[3]\ : CFG4
      generic map(INIT => x"0E00")

      port map(A => \fsmdet[5]_net_1\, B => \fsmdet[0]_net_1\, C
         => \SDAInt\, D => \SCLInt\, Y => N_861_i_0);
    
    \fsmsync_RNO[1]\ : CFG4
      generic map(INIT => x"3331")

      port map(A => N_995, B => \fsmsync_ns_i_1[6]_net_1\, C => 
        \fsmsync[1]_net_1\, D => \fsmsync[2]_net_1\, Y => 
        N_976_i_0);
    
    \fsmmod_ns_0[5]\ : CFG4
      generic map(INIT => x"FF40")

      port map(A => \SDAInt\, B => \fsmmod[6]_net_1\, C => 
        N_1059_1, D => N_1058, Y => \fsmmod_ns[5]\);
    
    \serSTA_WRITE_PROC.sersta_32_5[1]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \fsmsta[12]_net_1\, B => \fsmsta[24]_net_1\, 
        C => \COREI2C_0_2_INT[0]\, D => \fsmsta[28]_net_1\, Y => 
        \sersta_32_5[1]\);
    
    \serCON_WRITE_PROC.sercon_8_0_2[3]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \sercon[6]_net_1\, B => \COREI2C_0_2_INT[0]\, 
        C => \sercon_8_0_1[3]\, D => N_134, Y => 
        \sercon_8_0_2[3]\);
    
    \fsmsync[5]\ : SLE
      port map(D => N_968_i_0, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fsmsync[5]_net_1\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_i_m3[19]\ : CFG4
      generic map(INIT => x"F353")

      port map(A => \fsmsta[19]_net_1\, B => 
        \COREI2C_0_2_SDAO[0]\, C => N_2193, D => \un1_fsmsta_6\, 
        Y => N_2199);
    
    \serDAT_WRITE_PROC.serdat_9[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(2), B => 
        un105_ens1, C => \serdat[1]_net_1\, Y => \serdat_9[2]\);
    
    \FSMSYNC_SYNC_PROC.un141_ens1_2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \fsmsync[2]_net_1\, B => \fsmsync[5]_net_1\, 
        C => \fsmsync[6]_net_1\, D => \fsmsync[1]_net_1\, Y => 
        un141_ens1_2);
    
    \fsmmod_ns_i_0[2]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => \nedetect\, B => N_117_1, C => 
        \fsmmod[4]_net_1\, Y => \fsmmod_ns_i_0[2]_net_1\);
    
    \fsmmod_ns_i_o3_0_0[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREI2C_0_2_INT[0]\, B => \sercon[4]_net_1\, 
        Y => N_997);
    
    \sersta[2]\ : SLE
      port map(D => \sersta_32[2]\, CLK => FAB_CCC_GL0, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sersta[2]_net_1\);
    
    \CLK_COUNTER1_PROC.PCLK_count1_10[3]\ : CFG4
      generic map(INIT => x"060C")

      port map(A => \PCLK_count1[2]_net_1\, B => 
        \PCLK_count1[3]_net_1\, C => \un1_counter_rst_3\, D => 
        CO1, Y => \PCLK_count1_10[3]\);
    
    \FSMSTA_SYNC_PROC.fsmsta_8_ns_1[18]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => N_2181, B => un133_framesync, C => \ack\, D
         => un13_adrcompen, Y => \fsmsta_8_ns_1[18]\);
    
    un1_rtn_3 : CFG3
      generic map(INIT => x"81")

      port map(A => \SCLI_ff_reg[2]_net_1\, B => 
        \SCLI_ff_reg[1]_net_1\, C => \SCLI_ff_reg[0]_net_1\, Y
         => un1_rtn_3_1);
    
    nedetect_0_sqmuxa : CFG4
      generic map(INIT => x"0004")

      port map(A => \SCLI_ff_reg[0]_net_1\, B => \SCLInt\, C => 
        \SCLI_ff_reg[2]_net_1\, D => \SCLI_ff_reg[1]_net_1\, Y
         => \nedetect_0_sqmuxa\);
    
    starto_en_RNO : CFG3
      generic map(INIT => x"20")

      port map(A => \SCLInt\, B => \fsmmod[1]_net_1\, C => 
        \busfree\, Y => N_40_i_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREI2C_1 is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          COREI2C_0_2_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          MSS_READY                    : in    std_logic;
          FAB_CCC_GL0                  : in    std_logic;
          un3_penable                  : in    std_logic;
          bclke                        : in    std_logic;
          N_1218                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_2_SCL_IO_Y   : in    std_logic;
          BIBUF_COREI2C_0_2_SDA_IO_Y   : in    std_logic;
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un3_penable_1                : in    std_logic;
          un105_ens1_1                 : in    std_logic;
          N_40                         : in    std_logic;
          un5_penable_1                : in    std_logic
        );

end COREI2C_1;

architecture DEF_ARCH of COREI2C_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2CREAL_6_1
    port( COREI2C_0_2_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          seradr0apb                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          bclke                        : in    std_logic := 'U';
          N_1218                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_2_SCL_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_2_SDA_IO_Y   : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un3_penable_1                : in    std_logic := 'U';
          un105_ens1_1                 : in    std_logic := 'U';
          N_40                         : in    std_logic := 'U';
          un5_penable_1                : in    std_logic := 'U'
        );
  end component;

    signal \seradr0apb[4]_net_1\, VCC_net_1, GND_net_1, 
        \seradr0apb[5]_net_1\, \seradr0apb[6]_net_1\, 
        \seradr0apb[7]_net_1\, \seradr0apb[0]_net_1\, 
        \seradr0apb[1]_net_1\, \seradr0apb[2]_net_1\, 
        \seradr0apb[3]_net_1\ : std_logic;

    for all : COREI2CREAL_6_1
	Use entity work.COREI2CREAL_6_1(DEF_ARCH);
begin 


    \seradr0apb[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[7]_net_1\);
    
    \seradr0apb[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[6]_net_1\);
    
    \seradr0apb[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[2]_net_1\);
    
    \seradr0apb[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \seradr0apb[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[5]_net_1\);
    
    \seradr0apb[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[3]_net_1\);
    
    \seradr0apb[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[1]_net_1\);
    
    \seradr0apb[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        FAB_CCC_GL0, EN => un3_penable, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \seradr0apb[0]_net_1\);
    
    \G0a.0.ui2c\ : COREI2CREAL_6_1
      port map(COREI2C_0_2_SDAO_i(0) => COREI2C_0_2_SDAO_i(0), 
        COREI2C_0_2_SCLO_i(0) => COREI2C_0_2_SCLO_i(0), 
        COREI2C_0_2_INT(0) => COREI2C_0_2_INT(0), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), seradr0apb(7) => 
        \seradr0apb[7]_net_1\, seradr0apb(6) => 
        \seradr0apb[6]_net_1\, seradr0apb(5) => 
        \seradr0apb[5]_net_1\, seradr0apb(4) => 
        \seradr0apb[4]_net_1\, seradr0apb(3) => 
        \seradr0apb[3]_net_1\, seradr0apb(2) => 
        \seradr0apb[2]_net_1\, seradr0apb(1) => 
        \seradr0apb[1]_net_1\, seradr0apb(0) => 
        \seradr0apb[0]_net_1\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, bclke => bclke, N_1218 => 
        N_1218, N_1221 => N_1221, N_1217 => N_1217, N_1219 => 
        N_1219, N_1220 => N_1220, BIBUF_COREI2C_0_2_SCL_IO_Y => 
        BIBUF_COREI2C_0_2_SCL_IO_Y, BIBUF_COREI2C_0_2_SDA_IO_Y
         => BIBUF_COREI2C_0_2_SDA_IO_Y, N_1214 => N_1214, N_1215
         => N_1215, N_1216 => N_1216, un3_penable_1 => 
        un3_penable_1, un105_ens1_1 => un105_ens1_1, N_40 => N_40, 
        un5_penable_1 => un5_penable_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity M2sExt_sb is

    port( IO_0_Y             : in    std_logic_vector(0 to 0);
          GPIO_IN_c          : in    std_logic_vector(19 downto 4);
          GPIO_OUT_c         : out   std_logic_vector(2 downto 1);
          USB_ULPI_DATA      : inout std_logic_vector(7 downto 0) := (others => 'Z');
          COREI2C_0_6_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_6_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_5_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_5_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_4_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_4_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_3_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_3_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_2_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_2_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_1_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_1_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_0_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_0_SCL_IO : inout std_logic := 'Z';
          DEVRST_N           : in    std_logic;
          USB_RST_c          : out   std_logic;
          USB_ULPI_XCLK      : in    std_logic;
          USB_ULPI_STP       : out   std_logic;
          USB_ULPI_NXT       : in    std_logic;
          USB_ULPI_DIR       : in    std_logic
        );

end M2sExt_sb;

architecture DEF_ARCH of M2sExt_sb is 

  component M2sExt_sb_MSS
    port( USB_ULPI_DATA                               : inout   std_logic_vector(7 downto 0);
          GPOUT_reg                                   : in    std_logic_vector(3 to 3) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR  : inout   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                 : inout   std_logic_vector(8 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA                : out   std_logic_vector(31 downto 0);
          COREI2C_0_0_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_1_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_2_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_3_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_4_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_5_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          COREI2C_0_6_INT                             : in    std_logic_vector(0 to 0) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : in    std_logic_vector(31 downto 8) := (others => 'U');
          USB_ULPI_XCLK                               : in    std_logic := 'U';
          USB_ULPI_STP                                : out   std_logic;
          USB_ULPI_NXT                                : in    std_logic := 'U';
          USB_ULPI_DIR                                : in    std_logic := 'U';
          N_48                                        : in    std_logic := 'U';
          un561_psel_4                                : in    std_logic := 'U';
          m7_x                                        : in    std_logic := 'U';
          N_47                                        : in    std_logic := 'U';
          N_1217                                      : in    std_logic := 'U';
          N_1217_0                                    : in    std_logic := 'U';
          N_1217_1                                    : in    std_logic := 'U';
          N_1217_2                                    : in    std_logic := 'U';
          N_8_0                                       : in    std_logic := 'U';
          m71_1                                       : in    std_logic := 'U';
          N_1217_3                                    : in    std_logic := 'U';
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : inout   std_logic;
          CoreAPB3_0_APBmslave7_PSELx                 : in    std_logic := 'U';
          un30_psel                                   : in    std_logic := 'U';
          N_6186                                      : in    std_logic := 'U';
          M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N    : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE               : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                : out   std_logic;
          M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F         : out   std_logic;
          N_23_0_i_0                                  : in    std_logic := 'U';
          N_38_i_0                                    : in    std_logic := 'U';
          N_62_i_0                                    : in    std_logic := 'U';
          N_92_i_0                                    : in    std_logic := 'U';
          N_107_i_0                                   : in    std_logic := 'U';
          N_122_i_0                                   : in    std_logic := 'U';
          N_137_i_0                                   : in    std_logic := 'U';
          FAB_CCC_LOCK                                : in    std_logic := 'U';
          FAB_CCC_GL0                                 : in    std_logic := 'U'
        );
  end component;

  component COREI2C_2
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_3_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_3_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          un3_penable                  : in    std_logic := 'U';
          N_1217                       : out   std_logic;
          N_1218                       : out   std_logic;
          N_1220                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1221                       : out   std_logic;
          BIBUF_COREI2C_0_3_SDA_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_3_SCL_IO_Y   : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          bclke                        : in    std_logic := 'U';
          N_40                         : in    std_logic := 'U';
          un3_penable_1                : in    std_logic := 'U';
          un105_ens1_1                 : in    std_logic := 'U';
          un5_penable_1                : in    std_logic := 'U'
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CoreAPB3
    port( M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR  : in    std_logic_vector(15 downto 12) := (others => 'U');
          GPOUT_reg                                   : in    std_logic_vector(31 downto 20) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 8);
          CoreAPB3_0_APBmslave0_PADDR_8               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PADDR_7               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PADDR_0               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PADDR_6               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PADDR_5               : in    std_logic := 'U';
          INTR_reg_m_0                                : in    std_logic := 'U';
          INTR_reg_m_9                                : in    std_logic := 'U';
          INTR_reg_m_4                                : in    std_logic := 'U';
          INTR_reg_m_7                                : in    std_logic := 'U';
          INTR_reg_m_1                                : in    std_logic := 'U';
          N_8_0                                       : out   std_logic;
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : in    std_logic := 'U';
          m7_x                                        : out   std_logic;
          m46_1                                       : out   std_logic;
          N_122_i_1                                   : in    std_logic := 'U';
          N_122_i_0                                   : out   std_logic;
          N_92_i_1_1                                  : in    std_logic := 'U';
          N_92_i_0                                    : out   std_logic;
          N_48                                        : out   std_logic;
          m62_s                                       : in    std_logic := 'U';
          CONFIG_regror_28                            : in    std_logic := 'U';
          CONFIG_regror_29                            : in    std_logic := 'U';
          un561_psel_4                                : in    std_logic := 'U';
          N_1214                                      : in    std_logic := 'U';
          N_1215                                      : in    std_logic := 'U';
          N_1221                                      : in    std_logic := 'U';
          N_1219                                      : in    std_logic := 'U';
          N_1220                                      : in    std_logic := 'U';
          N_1218                                      : in    std_logic := 'U';
          N_1218_0                                    : in    std_logic := 'U';
          N_1218_1                                    : in    std_logic := 'U';
          N_1218_2                                    : in    std_logic := 'U';
          N_1216                                      : in    std_logic := 'U';
          N_1216_0                                    : in    std_logic := 'U';
          N_1216_1                                    : in    std_logic := 'U';
          N_1216_2                                    : in    std_logic := 'U';
          N_1216_3                                    : in    std_logic := 'U';
          N_1216_4                                    : in    std_logic := 'U';
          N_1214_0                                    : in    std_logic := 'U';
          N_1214_1                                    : in    std_logic := 'U';
          N_1214_2                                    : in    std_logic := 'U';
          N_1214_3                                    : in    std_logic := 'U';
          N_1214_4                                    : in    std_logic := 'U';
          N_1214_5                                    : in    std_logic := 'U';
          N_1217                                      : in    std_logic := 'U';
          N_1217_0                                    : in    std_logic := 'U';
          m71_1                                       : out   std_logic;
          N_1221_0                                    : in    std_logic := 'U';
          N_1221_1                                    : in    std_logic := 'U';
          N_1221_2                                    : in    std_logic := 'U';
          N_1221_3                                    : in    std_logic := 'U';
          N_1221_4                                    : in    std_logic := 'U';
          N_1221_5                                    : in    std_logic := 'U';
          N_1220_0                                    : in    std_logic := 'U';
          N_1220_1                                    : in    std_logic := 'U';
          N_1219_0                                    : in    std_logic := 'U';
          N_1219_1                                    : in    std_logic := 'U';
          N_1219_2                                    : in    std_logic := 'U';
          N_1219_3                                    : in    std_logic := 'U';
          N_1219_4                                    : in    std_logic := 'U';
          N_1219_5                                    : in    std_logic := 'U';
          N_1220_2                                    : in    std_logic := 'U';
          N_1220_3                                    : in    std_logic := 'U';
          N_1220_4                                    : in    std_logic := 'U';
          N_1220_5                                    : in    std_logic := 'U';
          N_1218_3                                    : in    std_logic := 'U';
          N_1218_4                                    : in    std_logic := 'U';
          N_1215_0                                    : in    std_logic := 'U';
          N_1215_1                                    : in    std_logic := 'U';
          N_1215_2                                    : in    std_logic := 'U';
          N_1215_3                                    : in    std_logic := 'U';
          N_1215_4                                    : in    std_logic := 'U';
          N_1215_5                                    : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE                : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE               : in    std_logic := 'U';
          CONFIG_rega23_1                             : in    std_logic := 'U';
          CoreAPB3_0_APBmslave7_PSELx                 : out   std_logic;
          N_1218_5                                    : in    std_logic := 'U';
          N_40                                        : out   std_logic;
          N_138                                       : out   std_logic;
          N_1216_5                                    : in    std_logic := 'U';
          N_43                                        : out   std_logic;
          un3_penable                                 : out   std_logic;
          un3_penable_0                               : out   std_logic;
          un3_penable_1                               : out   std_logic;
          un3_penable_2                               : out   std_logic;
          un3_penable_3                               : out   std_logic;
          un3_penable_4                               : out   std_logic;
          un3_penable_5                               : out   std_logic;
          N_24_0                                      : in    std_logic := 'U';
          N_137_i_0                                   : out   std_logic;
          N_37                                        : in    std_logic := 'U';
          N_107_i_0                                   : out   std_logic;
          N_53                                        : in    std_logic := 'U';
          N_62_i_0                                    : out   std_logic;
          N_58_0                                      : in    std_logic := 'U';
          N_38_i_0                                    : out   std_logic;
          N_63                                        : in    std_logic := 'U';
          N_23_0_i_0                                  : out   std_logic;
          N_440                                       : in    std_logic := 'U';
          un30_psel                                   : in    std_logic := 'U';
          N_438                                       : in    std_logic := 'U';
          N_439                                       : in    std_logic := 'U';
          N_435                                       : in    std_logic := 'U';
          N_441                                       : in    std_logic := 'U';
          N_437                                       : in    std_logic := 'U';
          N_436                                       : in    std_logic := 'U';
          N_338                                       : in    std_logic := 'U';
          N_333                                       : in    std_logic := 'U';
          N_310                                       : in    std_logic := 'U';
          N_419_mux                                   : in    std_logic := 'U';
          un3_prdata_o                                : in    std_logic := 'U';
          N_302                                       : in    std_logic := 'U';
          N_426_mux                                   : in    std_logic := 'U';
          N_345                                       : in    std_logic := 'U';
          N_421_mux                                   : in    std_logic := 'U';
          N_312                                       : in    std_logic := 'U';
          N_343                                       : in    std_logic := 'U';
          N_324                                       : in    std_logic := 'U';
          N_319                                       : in    std_logic := 'U';
          N_353                                       : in    std_logic := 'U';
          N_358                                       : in    std_logic := 'U';
          N_328                                       : in    std_logic := 'U'
        );
  end component;

  component CoreGPIO
    port( CoreAPB3_0_APBmslave0_PWDATA  : in    std_logic_vector(31 downto 0) := (others => 'U');
          GPIO_IN_c                     : in    std_logic_vector(19 downto 4) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR   : in    std_logic_vector(7 downto 0) := (others => 'U');
          GPIO_OUT_c                    : out   std_logic_vector(2 downto 1);
          GPOUT_reg_3                   : out   std_logic;
          GPOUT_reg_31                  : out   std_logic;
          GPOUT_reg_30                  : out   std_logic;
          GPOUT_reg_29                  : out   std_logic;
          GPOUT_reg_28                  : out   std_logic;
          GPOUT_reg_27                  : out   std_logic;
          GPOUT_reg_26                  : out   std_logic;
          GPOUT_reg_25                  : out   std_logic;
          GPOUT_reg_24                  : out   std_logic;
          GPOUT_reg_23                  : out   std_logic;
          GPOUT_reg_22                  : out   std_logic;
          GPOUT_reg_21                  : out   std_logic;
          GPOUT_reg_20                  : out   std_logic;
          INTR_reg_m_0                  : out   std_logic;
          INTR_reg_m_9                  : out   std_logic;
          INTR_reg_m_4                  : out   std_logic;
          INTR_reg_m_7                  : out   std_logic;
          INTR_reg_m_1                  : out   std_logic;
          MSS_READY                     : in    std_logic := 'U';
          FAB_CCC_GL0                   : in    std_logic := 'U';
          un30_psel                     : out   std_logic;
          m62_s                         : out   std_logic;
          un3_prdata_o                  : out   std_logic;
          CONFIG_regror_29              : out   std_logic;
          CONFIG_regror_28              : out   std_logic;
          N_24_0                        : out   std_logic;
          N_53                          : out   std_logic;
          N_58                          : out   std_logic;
          N_37                          : out   std_logic;
          N_122_i_1                     : out   std_logic;
          N_63                          : out   std_logic;
          N_92_i_1_1                    : out   std_logic;
          N_47                          : out   std_logic;
          N_310                         : out   std_logic;
          N_333                         : out   std_logic;
          N_338                         : out   std_logic;
          N_343                         : out   std_logic;
          N_319                         : out   std_logic;
          N_6186                        : out   std_logic;
          N_324                         : out   std_logic;
          N_353                         : out   std_logic;
          N_358                         : out   std_logic;
          N_328                         : out   std_logic;
          N_419_mux                     : out   std_logic;
          N_426_mux                     : out   std_logic;
          USB_RST_c                     : out   std_logic;
          N_421_mux                     : out   std_logic;
          CONFIG_rega23_1               : out   std_logic;
          CONFIG_rega20_2               : in    std_logic := 'U';
          N_48_1                        : in    std_logic := 'U';
          m46_1_0                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE  : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE : in    std_logic := 'U';
          CoreAPB3_0_APBmslave7_PSELx   : in    std_logic := 'U';
          N_438                         : out   std_logic;
          N_440                         : out   std_logic;
          N_439                         : out   std_logic;
          N_435                         : out   std_logic;
          N_441                         : out   std_logic;
          N_437                         : out   std_logic;
          N_436                         : out   std_logic;
          N_302                         : out   std_logic;
          N_345                         : out   std_logic;
          N_312                         : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREI2C
    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_0_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_0_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          un3_penable                                : in    std_logic := 'U';
          bclke                                      : out   std_logic;
          un561_psel_4                               : out   std_logic;
          CONFIG_rega20_2                            : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_0_SDA_IO_Y                 : in    std_logic := 'U';
          un105_ens1_3                               : out   std_logic;
          BIBUF_COREI2C_0_0_SCL_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          un3_penable_1                              : out   std_logic;
          un5_penable_0                              : out   std_logic;
          un105_ens1_0                               : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_138                                      : in    std_logic := 'U';
          un5_penable_2                              : in    std_logic := 'U'
        );
  end component;

  component CoreResetP
    port( MSS_READY                                : out   std_logic;
          FAB_CCC_GL0                              : in    std_logic := 'U';
          POWER_ON_RESET_N                         : in    std_logic := 'U';
          M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U'
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component COREI2C_0
    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_1_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_1_INT                            : out   std_logic_vector(0 to 0);
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(12 to 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(4 downto 0) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          un3_penable                                : in    std_logic := 'U';
          N_1221                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1218                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          BIBUF_COREI2C_0_1_SCL_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_1_SDA_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          un3_penable_1                              : out   std_logic;
          un105_ens1_3                               : in    std_logic := 'U';
          un105_ens1_1                               : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic := 'U';
          un5_penable_1                              : out   std_logic;
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          bclke                                      : in    std_logic := 'U';
          N_138                                      : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREI2C_4
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_5_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_5_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          un3_penable                  : in    std_logic := 'U';
          N_1218                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_5_SCL_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_5_SDA_IO_Y   : in    std_logic := 'U';
          bclke                        : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un105_ens1_0                 : in    std_logic := 'U';
          un105_ens1_3                 : in    std_logic := 'U';
          un3_penable_1                : in    std_logic := 'U';
          N_43                         : in    std_logic := 'U';
          un5_penable_0                : in    std_logic := 'U'
        );
  end component;

  component M2sExt_sb_CCC_0_FCCC
    port( IO_0_Y       : in    std_logic_vector(0 to 0) := (others => 'U');
          FAB_CCC_GL0  : out   std_logic;
          FAB_CCC_LOCK : out   std_logic
        );
  end component;

  component COREI2C_5
    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_6_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_6_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 2) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 12) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          un3_penable                                : in    std_logic := 'U';
          bclke                                      : in    std_logic := 'U';
          N_1218                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          BIBUF_COREI2C_0_6_SCL_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_6_SDA_IO_Y                 : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE              : in    std_logic := 'U';
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          N_8_0                                      : in    std_logic := 'U';
          un105_ens1_1                               : in    std_logic := 'U';
          un5_penable_1                              : in    std_logic := 'U'
        );
  end component;

  component COREI2C_3
    port( CoreAPB3_0_APBmslave0_PWDATA               : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_4_SDAO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_SCLO_i                         : out   std_logic_vector(0 to 0);
          COREI2C_0_4_INT                            : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR                : in    std_logic_vector(3 downto 1) := (others => 'U');
          M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(14 downto 13) := (others => 'U');
          MSS_READY                                  : in    std_logic := 'U';
          FAB_CCC_GL0                                : in    std_logic := 'U';
          un3_penable                                : in    std_logic := 'U';
          N_1218                                     : out   std_logic;
          N_1219                                     : out   std_logic;
          N_1217                                     : out   std_logic;
          N_1220                                     : out   std_logic;
          N_1221                                     : out   std_logic;
          BIBUF_COREI2C_0_4_SDA_IO_Y                 : in    std_logic := 'U';
          BIBUF_COREI2C_0_4_SCL_IO_Y                 : in    std_logic := 'U';
          N_1214                                     : out   std_logic;
          N_1215                                     : out   std_logic;
          N_1216                                     : out   std_logic;
          CONFIG_rega20_2                            : in    std_logic := 'U';
          un3_penable_1                              : in    std_logic := 'U';
          un105_ens1_3                               : in    std_logic := 'U';
          un5_penable_2                              : out   std_logic;
          bclke                                      : in    std_logic := 'U';
          N_8_0                                      : in    std_logic := 'U';
          N_43                                       : in    std_logic := 'U';
          un105_ens1_0                               : in    std_logic := 'U'
        );
  end component;

  component COREI2C_1
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREI2C_0_2_SDAO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_SCLO_i           : out   std_logic_vector(0 to 0);
          COREI2C_0_2_INT              : out   std_logic_vector(0 to 0);
          CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          MSS_READY                    : in    std_logic := 'U';
          FAB_CCC_GL0                  : in    std_logic := 'U';
          un3_penable                  : in    std_logic := 'U';
          bclke                        : in    std_logic := 'U';
          N_1218                       : out   std_logic;
          N_1221                       : out   std_logic;
          N_1217                       : out   std_logic;
          N_1219                       : out   std_logic;
          N_1220                       : out   std_logic;
          BIBUF_COREI2C_0_2_SCL_IO_Y   : in    std_logic := 'U';
          BIBUF_COREI2C_0_2_SDA_IO_Y   : in    std_logic := 'U';
          N_1214                       : out   std_logic;
          N_1215                       : out   std_logic;
          N_1216                       : out   std_logic;
          un3_penable_1                : in    std_logic := 'U';
          un105_ens1_1                 : in    std_logic := 'U';
          N_40                         : in    std_logic := 'U';
          un5_penable_1                : in    std_logic := 'U'
        );
  end component;

    signal BIBUF_COREI2C_0_6_SDA_IO_Y, GND_net_1, 
        \COREI2C_0_6_SDAO_i[0]\, BIBUF_COREI2C_0_6_SCL_IO_Y, 
        \COREI2C_0_6_SCLO_i[0]\, BIBUF_COREI2C_0_5_SDA_IO_Y, 
        \COREI2C_0_5_SDAO_i[0]\, BIBUF_COREI2C_0_5_SCL_IO_Y, 
        \COREI2C_0_5_SCLO_i[0]\, BIBUF_COREI2C_0_4_SDA_IO_Y, 
        \COREI2C_0_4_SDAO_i[0]\, BIBUF_COREI2C_0_4_SCL_IO_Y, 
        \COREI2C_0_4_SCLO_i[0]\, BIBUF_COREI2C_0_3_SDA_IO_Y, 
        \COREI2C_0_3_SDAO_i[0]\, BIBUF_COREI2C_0_3_SCL_IO_Y, 
        \COREI2C_0_3_SCLO_i[0]\, BIBUF_COREI2C_0_2_SDA_IO_Y, 
        \COREI2C_0_2_SDAO_i[0]\, BIBUF_COREI2C_0_2_SCL_IO_Y, 
        \COREI2C_0_2_SCLO_i[0]\, BIBUF_COREI2C_0_1_SDA_IO_Y, 
        \COREI2C_0_1_SDAO_i[0]\, BIBUF_COREI2C_0_1_SCL_IO_Y, 
        \COREI2C_0_1_SCLO_i[0]\, BIBUF_COREI2C_0_0_SDA_IO_Y, 
        \COREI2C_0_0_SDAO_i[0]\, BIBUF_COREI2C_0_0_SCL_IO_Y, 
        \COREI2C_0_0_SCLO_i[0]\, POWER_ON_RESET_N, FAB_CCC_GL0, 
        FAB_CCC_LOCK, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]\, 
        \CoreAPB3_0_APBmslave0_PADDR[8]\, 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, \GPOUT_reg[20]\, 
        \GPOUT_reg[21]\, \GPOUT_reg[22]\, \GPOUT_reg[23]\, 
        \GPOUT_reg[24]\, \GPOUT_reg[25]\, \GPOUT_reg[26]\, 
        \GPOUT_reg[27]\, \GPOUT_reg[28]\, \GPOUT_reg[29]\, 
        \GPOUT_reg[30]\, \GPOUT_reg[31]\, \INTR_reg_m[22]\, 
        \INTR_reg_m[31]\, \INTR_reg_m[26]\, \INTR_reg_m[29]\, 
        \INTR_reg_m[23]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\, 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\, N_8_0, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, m7_x, m46_1, 
        N_122_i_1, N_122_i_0, N_92_i_1_1, N_92_i_0, N_48, m62_s, 
        CONFIG_regror_28, CONFIG_regror_29, un561_psel_4, N_1214, 
        N_1215, N_1221, N_1219, N_1220, N_1218, N_1218_0, 
        N_1218_1, N_1218_2, N_1216, N_1216_0, N_1216_1, N_1216_2, 
        N_1216_3, N_1216_4, N_1214_0, N_1214_1, N_1214_2, 
        N_1214_3, N_1214_4, N_1214_5, N_1217, N_1217_0, m71_1, 
        N_1221_0, N_1221_1, N_1221_2, N_1221_3, N_1221_4, 
        N_1221_5, N_1220_0, N_1220_1, N_1219_0, N_1219_1, 
        N_1219_2, N_1219_3, N_1219_4, N_1219_5, N_1220_2, 
        N_1220_3, N_1220_4, N_1220_5, N_1218_3, N_1218_4, 
        N_1215_0, N_1215_1, N_1215_2, N_1215_3, N_1215_4, 
        N_1215_5, CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, CONFIG_rega23_1, 
        CoreAPB3_0_APBmslave7_PSELx, N_1218_5, N_40, N_138, 
        N_1216_5, N_43, un3_penable, un3_penable_0, un3_penable_1, 
        un3_penable_2, un3_penable_3, un3_penable_4, 
        un3_penable_5, N_24_0, N_137_i_0, N_37, N_107_i_0, N_53, 
        N_62_i_0, N_58, N_38_i_0, N_63, N_23_0_i_0, N_440, 
        un30_psel, N_438, N_439, N_435, N_441, N_437, N_436, 
        N_338, N_333, N_310, N_419_mux, un3_prdata_o, N_302, 
        N_426_mux, N_345, N_421_mux, N_312, N_343, N_324, N_319, 
        N_353, N_358, N_328, \GPOUT_reg[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[8]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[9]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[10]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[11]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[12]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[13]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[14]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[15]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[16]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[17]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[18]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[19]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[20]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[21]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[22]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[23]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[24]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[25]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[26]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[27]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[28]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[29]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[30]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[31]\, 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, MSS_READY, N_47, N_6186, 
        CONFIG_rega20_2, \COREI2C_0_0_INT[0]\, bclke, N_1217_1, 
        un105_ens1_3, un3_penable_1_0, un5_penable_0, 
        un105_ens1_0, un5_penable_2, \COREI2C_0_1_INT[0]\, 
        un3_penable_1_1, un105_ens1_1, un5_penable_1, 
        \COREI2C_0_2_INT[0]\, N_1217_2, \COREI2C_0_3_INT[0]\, 
        N_1217_3, \COREI2C_0_4_INT[0]\, N_1217_4, 
        \COREI2C_0_5_INT[0]\, \COREI2C_0_6_INT[0]\, N_1217_5, 
        M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, VCC_net_1
         : std_logic;

    for all : M2sExt_sb_MSS
	Use entity work.M2sExt_sb_MSS(DEF_ARCH);
    for all : COREI2C_2
	Use entity work.COREI2C_2(DEF_ARCH);
    for all : CoreAPB3
	Use entity work.CoreAPB3(DEF_ARCH);
    for all : CoreGPIO
	Use entity work.CoreGPIO(DEF_ARCH);
    for all : COREI2C
	Use entity work.COREI2C(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : COREI2C_0
	Use entity work.COREI2C_0(DEF_ARCH);
    for all : COREI2C_4
	Use entity work.COREI2C_4(DEF_ARCH);
    for all : M2sExt_sb_CCC_0_FCCC
	Use entity work.M2sExt_sb_CCC_0_FCCC(DEF_ARCH);
    for all : COREI2C_5
	Use entity work.COREI2C_5(DEF_ARCH);
    for all : COREI2C_3
	Use entity work.COREI2C_3(DEF_ARCH);
    for all : COREI2C_1
	Use entity work.COREI2C_1(DEF_ARCH);
begin 


    M2sExt_sb_MSS_0 : M2sExt_sb_MSS
      port map(USB_ULPI_DATA(7) => USB_ULPI_DATA(7), 
        USB_ULPI_DATA(6) => USB_ULPI_DATA(6), USB_ULPI_DATA(5)
         => USB_ULPI_DATA(5), USB_ULPI_DATA(4) => 
        USB_ULPI_DATA(4), USB_ULPI_DATA(3) => USB_ULPI_DATA(3), 
        USB_ULPI_DATA(2) => USB_ULPI_DATA(2), USB_ULPI_DATA(1)
         => USB_ULPI_DATA(1), USB_ULPI_DATA(0) => 
        USB_ULPI_DATA(0), GPOUT_reg(3) => \GPOUT_reg[3]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PADDR(8) => 
        \CoreAPB3_0_APBmslave0_PADDR[8]\, 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(31) => 
        \CoreAPB3_0_APBmslave0_PWDATA[31]\, 
        CoreAPB3_0_APBmslave0_PWDATA(30) => 
        \CoreAPB3_0_APBmslave0_PWDATA[30]\, 
        CoreAPB3_0_APBmslave0_PWDATA(29) => 
        \CoreAPB3_0_APBmslave0_PWDATA[29]\, 
        CoreAPB3_0_APBmslave0_PWDATA(28) => 
        \CoreAPB3_0_APBmslave0_PWDATA[28]\, 
        CoreAPB3_0_APBmslave0_PWDATA(27) => 
        \CoreAPB3_0_APBmslave0_PWDATA[27]\, 
        CoreAPB3_0_APBmslave0_PWDATA(26) => 
        \CoreAPB3_0_APBmslave0_PWDATA[26]\, 
        CoreAPB3_0_APBmslave0_PWDATA(25) => 
        \CoreAPB3_0_APBmslave0_PWDATA[25]\, 
        CoreAPB3_0_APBmslave0_PWDATA(24) => 
        \CoreAPB3_0_APBmslave0_PWDATA[24]\, 
        CoreAPB3_0_APBmslave0_PWDATA(23) => 
        \CoreAPB3_0_APBmslave0_PWDATA[23]\, 
        CoreAPB3_0_APBmslave0_PWDATA(22) => 
        \CoreAPB3_0_APBmslave0_PWDATA[22]\, 
        CoreAPB3_0_APBmslave0_PWDATA(21) => 
        \CoreAPB3_0_APBmslave0_PWDATA[21]\, 
        CoreAPB3_0_APBmslave0_PWDATA(20) => 
        \CoreAPB3_0_APBmslave0_PWDATA[20]\, 
        CoreAPB3_0_APBmslave0_PWDATA(19) => 
        \CoreAPB3_0_APBmslave0_PWDATA[19]\, 
        CoreAPB3_0_APBmslave0_PWDATA(18) => 
        \CoreAPB3_0_APBmslave0_PWDATA[18]\, 
        CoreAPB3_0_APBmslave0_PWDATA(17) => 
        \CoreAPB3_0_APBmslave0_PWDATA[17]\, 
        CoreAPB3_0_APBmslave0_PWDATA(16) => 
        \CoreAPB3_0_APBmslave0_PWDATA[16]\, 
        CoreAPB3_0_APBmslave0_PWDATA(15) => 
        \CoreAPB3_0_APBmslave0_PWDATA[15]\, 
        CoreAPB3_0_APBmslave0_PWDATA(14) => 
        \CoreAPB3_0_APBmslave0_PWDATA[14]\, 
        CoreAPB3_0_APBmslave0_PWDATA(13) => 
        \CoreAPB3_0_APBmslave0_PWDATA[13]\, 
        CoreAPB3_0_APBmslave0_PWDATA(12) => 
        \CoreAPB3_0_APBmslave0_PWDATA[12]\, 
        CoreAPB3_0_APBmslave0_PWDATA(11) => 
        \CoreAPB3_0_APBmslave0_PWDATA[11]\, 
        CoreAPB3_0_APBmslave0_PWDATA(10) => 
        \CoreAPB3_0_APBmslave0_PWDATA[10]\, 
        CoreAPB3_0_APBmslave0_PWDATA(9) => 
        \CoreAPB3_0_APBmslave0_PWDATA[9]\, 
        CoreAPB3_0_APBmslave0_PWDATA(8) => 
        \CoreAPB3_0_APBmslave0_PWDATA[8]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_0_INT(0) => 
        \COREI2C_0_0_INT[0]\, COREI2C_0_1_INT(0) => 
        \COREI2C_0_1_INT[0]\, COREI2C_0_2_INT(0) => 
        \COREI2C_0_2_INT[0]\, COREI2C_0_3_INT(0) => 
        \COREI2C_0_3_INT[0]\, COREI2C_0_4_INT(0) => 
        \COREI2C_0_4_INT[0]\, COREI2C_0_5_INT(0) => 
        \COREI2C_0_5_INT[0]\, COREI2C_0_6_INT(0) => 
        \COREI2C_0_6_INT[0]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\, 
        USB_ULPI_XCLK => USB_ULPI_XCLK, USB_ULPI_STP => 
        USB_ULPI_STP, USB_ULPI_NXT => USB_ULPI_NXT, USB_ULPI_DIR
         => USB_ULPI_DIR, N_48 => N_48, un561_psel_4 => 
        un561_psel_4, m7_x => m7_x, N_47 => N_47, N_1217 => 
        N_1217_5, N_1217_0 => N_1217_4, N_1217_1 => N_1217_1, 
        N_1217_2 => N_1217_2, N_8_0 => N_8_0, m71_1 => m71_1, 
        N_1217_3 => N_1217_3, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave7_PSELx => 
        CoreAPB3_0_APBmslave7_PSELx, un30_psel => un30_psel, 
        N_6186 => N_6186, 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, N_23_0_i_0 => 
        N_23_0_i_0, N_38_i_0 => N_38_i_0, N_62_i_0 => N_62_i_0, 
        N_92_i_0 => N_92_i_0, N_107_i_0 => N_107_i_0, N_122_i_0
         => N_122_i_0, N_137_i_0 => N_137_i_0, FAB_CCC_LOCK => 
        FAB_CCC_LOCK, FAB_CCC_GL0 => FAB_CCC_GL0);
    
    COREI2C_0_3 : COREI2C_2
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_3_SDAO_i(0)
         => \COREI2C_0_3_SDAO_i[0]\, COREI2C_0_3_SCLO_i(0) => 
        \COREI2C_0_3_SCLO_i[0]\, COREI2C_0_3_INT(0) => 
        \COREI2C_0_3_INT[0]\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, un3_penable => un3_penable_5, 
        N_1217 => N_1217_3, N_1218 => N_1218_5, N_1220 => N_1220, 
        N_1219 => N_1219, N_1221 => N_1221, 
        BIBUF_COREI2C_0_3_SDA_IO_Y => BIBUF_COREI2C_0_3_SDA_IO_Y, 
        BIBUF_COREI2C_0_3_SCL_IO_Y => BIBUF_COREI2C_0_3_SCL_IO_Y, 
        N_1214 => N_1214, N_1215 => N_1215, N_1216 => N_1216_5, 
        bclke => bclke, N_40 => N_40, un3_penable_1 => 
        un3_penable_1_1, un105_ens1_1 => un105_ens1_1, 
        un5_penable_1 => un5_penable_1);
    
    BIBUF_COREI2C_0_3_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_3_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_3_SCLO_i[0]\, Y => BIBUF_COREI2C_0_3_SCL_IO_Y);
    
    CoreAPB3_0 : CoreAPB3
      port map(M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(15) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        GPOUT_reg(31) => \GPOUT_reg[31]\, GPOUT_reg(30) => 
        \GPOUT_reg[30]\, GPOUT_reg(29) => \GPOUT_reg[29]\, 
        GPOUT_reg(28) => \GPOUT_reg[28]\, GPOUT_reg(27) => 
        \GPOUT_reg[27]\, GPOUT_reg(26) => \GPOUT_reg[26]\, 
        GPOUT_reg(25) => \GPOUT_reg[25]\, GPOUT_reg(24) => 
        \GPOUT_reg[24]\, GPOUT_reg(23) => \GPOUT_reg[23]\, 
        GPOUT_reg(22) => \GPOUT_reg[22]\, GPOUT_reg(21) => 
        \GPOUT_reg[21]\, GPOUT_reg(20) => \GPOUT_reg[20]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\, 
        CoreAPB3_0_APBmslave0_PADDR_8 => 
        \CoreAPB3_0_APBmslave0_PADDR[8]\, 
        CoreAPB3_0_APBmslave0_PADDR_7 => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR_0 => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        CoreAPB3_0_APBmslave0_PADDR_6 => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR_5 => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, INTR_reg_m_0 => 
        \INTR_reg_m[22]\, INTR_reg_m_9 => \INTR_reg_m[31]\, 
        INTR_reg_m_4 => \INTR_reg_m[26]\, INTR_reg_m_7 => 
        \INTR_reg_m[29]\, INTR_reg_m_1 => \INTR_reg_m[23]\, N_8_0
         => N_8_0, M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx => 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, m7_x => m7_x, 
        m46_1 => m46_1, N_122_i_1 => N_122_i_1, N_122_i_0 => 
        N_122_i_0, N_92_i_1_1 => N_92_i_1_1, N_92_i_0 => N_92_i_0, 
        N_48 => N_48, m62_s => m62_s, CONFIG_regror_28 => 
        CONFIG_regror_28, CONFIG_regror_29 => CONFIG_regror_29, 
        un561_psel_4 => un561_psel_4, N_1214 => N_1214, N_1215
         => N_1215, N_1221 => N_1221, N_1219 => N_1219, N_1220
         => N_1220, N_1218 => N_1218, N_1218_0 => N_1218_0, 
        N_1218_1 => N_1218_1, N_1218_2 => N_1218_2, N_1216 => 
        N_1216, N_1216_0 => N_1216_0, N_1216_1 => N_1216_1, 
        N_1216_2 => N_1216_2, N_1216_3 => N_1216_3, N_1216_4 => 
        N_1216_4, N_1214_0 => N_1214_0, N_1214_1 => N_1214_1, 
        N_1214_2 => N_1214_2, N_1214_3 => N_1214_3, N_1214_4 => 
        N_1214_4, N_1214_5 => N_1214_5, N_1217 => N_1217, 
        N_1217_0 => N_1217_0, m71_1 => m71_1, N_1221_0 => 
        N_1221_0, N_1221_1 => N_1221_1, N_1221_2 => N_1221_2, 
        N_1221_3 => N_1221_3, N_1221_4 => N_1221_4, N_1221_5 => 
        N_1221_5, N_1220_0 => N_1220_0, N_1220_1 => N_1220_1, 
        N_1219_0 => N_1219_0, N_1219_1 => N_1219_1, N_1219_2 => 
        N_1219_2, N_1219_3 => N_1219_3, N_1219_4 => N_1219_4, 
        N_1219_5 => N_1219_5, N_1220_2 => N_1220_2, N_1220_3 => 
        N_1220_3, N_1220_4 => N_1220_4, N_1220_5 => N_1220_5, 
        N_1218_3 => N_1218_3, N_1218_4 => N_1218_4, N_1215_0 => 
        N_1215_0, N_1215_1 => N_1215_1, N_1215_2 => N_1215_2, 
        N_1215_3 => N_1215_3, N_1215_4 => N_1215_4, N_1215_5 => 
        N_1215_5, CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, CONFIG_rega23_1 => 
        CONFIG_rega23_1, CoreAPB3_0_APBmslave7_PSELx => 
        CoreAPB3_0_APBmslave7_PSELx, N_1218_5 => N_1218_5, N_40
         => N_40, N_138 => N_138, N_1216_5 => N_1216_5, N_43 => 
        N_43, un3_penable => un3_penable, un3_penable_0 => 
        un3_penable_0, un3_penable_1 => un3_penable_1, 
        un3_penable_2 => un3_penable_2, un3_penable_3 => 
        un3_penable_3, un3_penable_4 => un3_penable_4, 
        un3_penable_5 => un3_penable_5, N_24_0 => N_24_0, 
        N_137_i_0 => N_137_i_0, N_37 => N_37, N_107_i_0 => 
        N_107_i_0, N_53 => N_53, N_62_i_0 => N_62_i_0, N_58_0 => 
        N_58, N_38_i_0 => N_38_i_0, N_63 => N_63, N_23_0_i_0 => 
        N_23_0_i_0, N_440 => N_440, un30_psel => un30_psel, N_438
         => N_438, N_439 => N_439, N_435 => N_435, N_441 => N_441, 
        N_437 => N_437, N_436 => N_436, N_338 => N_338, N_333 => 
        N_333, N_310 => N_310, N_419_mux => N_419_mux, 
        un3_prdata_o => un3_prdata_o, N_302 => N_302, N_426_mux
         => N_426_mux, N_345 => N_345, N_421_mux => N_421_mux, 
        N_312 => N_312, N_343 => N_343, N_324 => N_324, N_319 => 
        N_319, N_353 => N_353, N_358 => N_358, N_328 => N_328);
    
    BIBUF_COREI2C_0_6_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_6_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_6_SCLO_i[0]\, Y => BIBUF_COREI2C_0_6_SCL_IO_Y);
    
    BIBUF_COREI2C_0_4_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_4_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_4_SCLO_i[0]\, Y => BIBUF_COREI2C_0_4_SCL_IO_Y);
    
    BIBUF_COREI2C_0_0_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_0_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_0_SDAO_i[0]\, Y => BIBUF_COREI2C_0_0_SDA_IO_Y);
    
    CoreGPIO_0_0 : CoreGPIO
      port map(CoreAPB3_0_APBmslave0_PWDATA(31) => 
        \CoreAPB3_0_APBmslave0_PWDATA[31]\, 
        CoreAPB3_0_APBmslave0_PWDATA(30) => 
        \CoreAPB3_0_APBmslave0_PWDATA[30]\, 
        CoreAPB3_0_APBmslave0_PWDATA(29) => 
        \CoreAPB3_0_APBmslave0_PWDATA[29]\, 
        CoreAPB3_0_APBmslave0_PWDATA(28) => 
        \CoreAPB3_0_APBmslave0_PWDATA[28]\, 
        CoreAPB3_0_APBmslave0_PWDATA(27) => 
        \CoreAPB3_0_APBmslave0_PWDATA[27]\, 
        CoreAPB3_0_APBmslave0_PWDATA(26) => 
        \CoreAPB3_0_APBmslave0_PWDATA[26]\, 
        CoreAPB3_0_APBmslave0_PWDATA(25) => 
        \CoreAPB3_0_APBmslave0_PWDATA[25]\, 
        CoreAPB3_0_APBmslave0_PWDATA(24) => 
        \CoreAPB3_0_APBmslave0_PWDATA[24]\, 
        CoreAPB3_0_APBmslave0_PWDATA(23) => 
        \CoreAPB3_0_APBmslave0_PWDATA[23]\, 
        CoreAPB3_0_APBmslave0_PWDATA(22) => 
        \CoreAPB3_0_APBmslave0_PWDATA[22]\, 
        CoreAPB3_0_APBmslave0_PWDATA(21) => 
        \CoreAPB3_0_APBmslave0_PWDATA[21]\, 
        CoreAPB3_0_APBmslave0_PWDATA(20) => 
        \CoreAPB3_0_APBmslave0_PWDATA[20]\, 
        CoreAPB3_0_APBmslave0_PWDATA(19) => 
        \CoreAPB3_0_APBmslave0_PWDATA[19]\, 
        CoreAPB3_0_APBmslave0_PWDATA(18) => 
        \CoreAPB3_0_APBmslave0_PWDATA[18]\, 
        CoreAPB3_0_APBmslave0_PWDATA(17) => 
        \CoreAPB3_0_APBmslave0_PWDATA[17]\, 
        CoreAPB3_0_APBmslave0_PWDATA(16) => 
        \CoreAPB3_0_APBmslave0_PWDATA[16]\, 
        CoreAPB3_0_APBmslave0_PWDATA(15) => 
        \CoreAPB3_0_APBmslave0_PWDATA[15]\, 
        CoreAPB3_0_APBmslave0_PWDATA(14) => 
        \CoreAPB3_0_APBmslave0_PWDATA[14]\, 
        CoreAPB3_0_APBmslave0_PWDATA(13) => 
        \CoreAPB3_0_APBmslave0_PWDATA[13]\, 
        CoreAPB3_0_APBmslave0_PWDATA(12) => 
        \CoreAPB3_0_APBmslave0_PWDATA[12]\, 
        CoreAPB3_0_APBmslave0_PWDATA(11) => 
        \CoreAPB3_0_APBmslave0_PWDATA[11]\, 
        CoreAPB3_0_APBmslave0_PWDATA(10) => 
        \CoreAPB3_0_APBmslave0_PWDATA[10]\, 
        CoreAPB3_0_APBmslave0_PWDATA(9) => 
        \CoreAPB3_0_APBmslave0_PWDATA[9]\, 
        CoreAPB3_0_APBmslave0_PWDATA(8) => 
        \CoreAPB3_0_APBmslave0_PWDATA[8]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, GPIO_IN_c(19) => 
        GPIO_IN_c(19), GPIO_IN_c(18) => GPIO_IN_c(18), 
        GPIO_IN_c(17) => GPIO_IN_c(17), GPIO_IN_c(16) => 
        GPIO_IN_c(16), GPIO_IN_c(15) => GPIO_IN_c(15), 
        GPIO_IN_c(14) => GPIO_IN_c(14), GPIO_IN_c(13) => 
        GPIO_IN_c(13), GPIO_IN_c(12) => GPIO_IN_c(12), 
        GPIO_IN_c(11) => GPIO_IN_c(11), GPIO_IN_c(10) => 
        GPIO_IN_c(10), GPIO_IN_c(9) => GPIO_IN_c(9), GPIO_IN_c(8)
         => GPIO_IN_c(8), GPIO_IN_c(7) => GPIO_IN_c(7), 
        GPIO_IN_c(6) => GPIO_IN_c(6), GPIO_IN_c(5) => 
        GPIO_IN_c(5), GPIO_IN_c(4) => GPIO_IN_c(4), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, GPIO_OUT_c(2) => 
        GPIO_OUT_c(2), GPIO_OUT_c(1) => GPIO_OUT_c(1), 
        GPOUT_reg_3 => \GPOUT_reg[3]\, GPOUT_reg_31 => 
        \GPOUT_reg[31]\, GPOUT_reg_30 => \GPOUT_reg[30]\, 
        GPOUT_reg_29 => \GPOUT_reg[29]\, GPOUT_reg_28 => 
        \GPOUT_reg[28]\, GPOUT_reg_27 => \GPOUT_reg[27]\, 
        GPOUT_reg_26 => \GPOUT_reg[26]\, GPOUT_reg_25 => 
        \GPOUT_reg[25]\, GPOUT_reg_24 => \GPOUT_reg[24]\, 
        GPOUT_reg_23 => \GPOUT_reg[23]\, GPOUT_reg_22 => 
        \GPOUT_reg[22]\, GPOUT_reg_21 => \GPOUT_reg[21]\, 
        GPOUT_reg_20 => \GPOUT_reg[20]\, INTR_reg_m_0 => 
        \INTR_reg_m[22]\, INTR_reg_m_9 => \INTR_reg_m[31]\, 
        INTR_reg_m_4 => \INTR_reg_m[26]\, INTR_reg_m_7 => 
        \INTR_reg_m[29]\, INTR_reg_m_1 => \INTR_reg_m[23]\, 
        MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        un30_psel => un30_psel, m62_s => m62_s, un3_prdata_o => 
        un3_prdata_o, CONFIG_regror_29 => CONFIG_regror_29, 
        CONFIG_regror_28 => CONFIG_regror_28, N_24_0 => N_24_0, 
        N_53 => N_53, N_58 => N_58, N_37 => N_37, N_122_i_1 => 
        N_122_i_1, N_63 => N_63, N_92_i_1_1 => N_92_i_1_1, N_47
         => N_47, N_310 => N_310, N_333 => N_333, N_338 => N_338, 
        N_343 => N_343, N_319 => N_319, N_6186 => N_6186, N_324
         => N_324, N_353 => N_353, N_358 => N_358, N_328 => N_328, 
        N_419_mux => N_419_mux, N_426_mux => N_426_mux, USB_RST_c
         => USB_RST_c, N_421_mux => N_421_mux, CONFIG_rega23_1
         => CONFIG_rega23_1, CONFIG_rega20_2 => CONFIG_rega20_2, 
        N_48_1 => N_48, m46_1_0 => m46_1, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave7_PSELx => 
        CoreAPB3_0_APBmslave7_PSELx, N_438 => N_438, N_440 => 
        N_440, N_439 => N_439, N_435 => N_435, N_441 => N_441, 
        N_437 => N_437, N_436 => N_436, N_302 => N_302, N_345 => 
        N_345, N_312 => N_312);
    
    BIBUF_COREI2C_0_2_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_2_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_2_SDAO_i[0]\, Y => BIBUF_COREI2C_0_2_SDA_IO_Y);
    
    BIBUF_COREI2C_0_1_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_1_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_1_SCLO_i[0]\, Y => BIBUF_COREI2C_0_1_SCL_IO_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    COREI2C_0_0 : COREI2C
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_0_SDAO_i(0)
         => \COREI2C_0_0_SDAO_i[0]\, COREI2C_0_0_SCLO_i(0) => 
        \COREI2C_0_0_SCLO_i[0]\, COREI2C_0_0_INT(0) => 
        \COREI2C_0_0_INT[0]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, un3_penable => un3_penable_3, 
        bclke => bclke, un561_psel_4 => un561_psel_4, 
        CONFIG_rega20_2 => CONFIG_rega20_2, N_1221 => N_1221_1, 
        N_1217 => N_1217_1, N_1220 => N_1220_3, N_1218 => 
        N_1218_0, N_1219 => N_1219_3, BIBUF_COREI2C_0_0_SDA_IO_Y
         => BIBUF_COREI2C_0_0_SDA_IO_Y, un105_ens1_3 => 
        un105_ens1_3, BIBUF_COREI2C_0_0_SCL_IO_Y => 
        BIBUF_COREI2C_0_0_SCL_IO_Y, CoreAPB3_0_APBmslave0_PENABLE
         => CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, un3_penable_1 => 
        un3_penable_1_0, un5_penable_0 => un5_penable_0, 
        un105_ens1_0 => un105_ens1_0, N_1214 => N_1214_5, N_1215
         => N_1215_1, N_1216 => N_1216_0, N_138 => N_138, 
        un5_penable_2 => un5_penable_2);
    
    BIBUF_COREI2C_0_6_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_6_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_6_SDAO_i[0]\, Y => BIBUF_COREI2C_0_6_SDA_IO_Y);
    
    CORERESETP_0 : CoreResetP
      port map(MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        POWER_ON_RESET_N => POWER_ON_RESET_N, 
        M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        M2sExt_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        M2sExt_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => POWER_ON_RESET_N, DEVRST_N => 
        DEVRST_N);
    
    BIBUF_COREI2C_0_3_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_3_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_3_SDAO_i[0]\, Y => BIBUF_COREI2C_0_3_SDA_IO_Y);
    
    COREI2C_0_1 : COREI2C_0
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_1_SDAO_i(0)
         => \COREI2C_0_1_SDAO_i[0]\, COREI2C_0_1_SCLO_i(0) => 
        \COREI2C_0_1_SCLO_i[0]\, COREI2C_0_1_INT(0) => 
        \COREI2C_0_1_INT[0]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, un3_penable => un3_penable_2, 
        N_1221 => N_1221_5, N_1217 => N_1217_0, N_1218 => 
        N_1218_4, N_1220 => N_1220_1, N_1219 => N_1219_1, 
        BIBUF_COREI2C_0_1_SCL_IO_Y => BIBUF_COREI2C_0_1_SCL_IO_Y, 
        BIBUF_COREI2C_0_1_SDA_IO_Y => BIBUF_COREI2C_0_1_SDA_IO_Y, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, un3_penable_1 => 
        un3_penable_1_1, un105_ens1_3 => un105_ens1_3, 
        un105_ens1_1 => un105_ens1_1, CONFIG_rega20_2 => 
        CONFIG_rega20_2, un5_penable_1 => un5_penable_1, N_1214
         => N_1214_1, N_1215 => N_1215_5, N_1216 => N_1216_4, 
        bclke => bclke, N_138 => N_138);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    BIBUF_COREI2C_0_2_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_2_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_2_SCLO_i[0]\, Y => BIBUF_COREI2C_0_2_SCL_IO_Y);
    
    COREI2C_0_5 : COREI2C_4
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_5_SDAO_i(0)
         => \COREI2C_0_5_SDAO_i[0]\, COREI2C_0_5_SCLO_i(0) => 
        \COREI2C_0_5_SCLO_i[0]\, COREI2C_0_5_INT(0) => 
        \COREI2C_0_5_INT[0]\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, un3_penable => un3_penable_0, 
        N_1218 => N_1218_3, N_1217 => N_1217, N_1221 => N_1221_4, 
        N_1219 => N_1219_0, N_1220 => N_1220_0, 
        BIBUF_COREI2C_0_5_SCL_IO_Y => BIBUF_COREI2C_0_5_SCL_IO_Y, 
        BIBUF_COREI2C_0_5_SDA_IO_Y => BIBUF_COREI2C_0_5_SDA_IO_Y, 
        bclke => bclke, N_1214 => N_1214_0, N_1215 => N_1215_4, 
        N_1216 => N_1216_3, un105_ens1_0 => un105_ens1_0, 
        un105_ens1_3 => un105_ens1_3, un3_penable_1 => 
        un3_penable_1_1, N_43 => N_43, un5_penable_0 => 
        un5_penable_0);
    
    CCC_0 : M2sExt_sb_CCC_0_FCCC
      port map(IO_0_Y(0) => IO_0_Y(0), FAB_CCC_GL0 => FAB_CCC_GL0, 
        FAB_CCC_LOCK => FAB_CCC_LOCK);
    
    BIBUF_COREI2C_0_0_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_0_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_0_SCLO_i[0]\, Y => BIBUF_COREI2C_0_0_SCL_IO_Y);
    
    BIBUF_COREI2C_0_5_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_5_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_5_SDAO_i[0]\, Y => BIBUF_COREI2C_0_5_SDA_IO_Y);
    
    BIBUF_COREI2C_0_5_SCL_IO : BIBUF
      port map(PAD => COREI2C_0_5_SCL_IO, D => GND_net_1, E => 
        \COREI2C_0_5_SCLO_i[0]\, Y => BIBUF_COREI2C_0_5_SCL_IO_Y);
    
    COREI2C_0_6 : COREI2C_5
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_6_SDAO_i(0)
         => \COREI2C_0_6_SDAO_i[0]\, COREI2C_0_6_SCLO_i(0) => 
        \COREI2C_0_6_SCLO_i[0]\, COREI2C_0_6_INT(0) => 
        \COREI2C_0_6_INT[0]\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(12) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]\, 
        MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        un3_penable => un3_penable, bclke => bclke, N_1218 => 
        N_1218_1, N_1221 => N_1221_2, N_1219 => N_1219_4, N_1217
         => N_1217_5, N_1220 => N_1220_4, 
        BIBUF_COREI2C_0_6_SCL_IO_Y => BIBUF_COREI2C_0_6_SCL_IO_Y, 
        BIBUF_COREI2C_0_6_SDA_IO_Y => BIBUF_COREI2C_0_6_SDA_IO_Y, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, N_1214 => N_1214_2, N_1215
         => N_1215_2, N_1216 => N_1216_1, N_8_0 => N_8_0, 
        un105_ens1_1 => un105_ens1_1, un5_penable_1 => 
        un5_penable_1);
    
    COREI2C_0_4 : COREI2C_3
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_4_SDAO_i(0)
         => \COREI2C_0_4_SDAO_i[0]\, COREI2C_0_4_SCLO_i(0) => 
        \COREI2C_0_4_SCLO_i[0]\, COREI2C_0_4_INT(0) => 
        \COREI2C_0_4_INT[0]\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(14) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]\, 
        M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR(13) => 
        \M2sExt_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]\, 
        MSS_READY => MSS_READY, FAB_CCC_GL0 => FAB_CCC_GL0, 
        un3_penable => un3_penable_1, N_1218 => N_1218, N_1219
         => N_1219_2, N_1217 => N_1217_4, N_1220 => N_1220_2, 
        N_1221 => N_1221_0, BIBUF_COREI2C_0_4_SDA_IO_Y => 
        BIBUF_COREI2C_0_4_SDA_IO_Y, BIBUF_COREI2C_0_4_SCL_IO_Y
         => BIBUF_COREI2C_0_4_SCL_IO_Y, N_1214 => N_1214_4, 
        N_1215 => N_1215_0, N_1216 => N_1216, CONFIG_rega20_2 => 
        CONFIG_rega20_2, un3_penable_1 => un3_penable_1_0, 
        un105_ens1_3 => un105_ens1_3, un5_penable_2 => 
        un5_penable_2, bclke => bclke, N_8_0 => N_8_0, N_43 => 
        N_43, un105_ens1_0 => un105_ens1_0);
    
    BIBUF_COREI2C_0_1_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_1_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_1_SDAO_i[0]\, Y => BIBUF_COREI2C_0_1_SDA_IO_Y);
    
    COREI2C_0_2 : COREI2C_1
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, COREI2C_0_2_SDAO_i(0)
         => \COREI2C_0_2_SDAO_i[0]\, COREI2C_0_2_SCLO_i(0) => 
        \COREI2C_0_2_SCLO_i[0]\, COREI2C_0_2_INT(0) => 
        \COREI2C_0_2_INT[0]\, CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, MSS_READY => MSS_READY, 
        FAB_CCC_GL0 => FAB_CCC_GL0, un3_penable => un3_penable_4, 
        bclke => bclke, N_1218 => N_1218_2, N_1221 => N_1221_3, 
        N_1217 => N_1217_2, N_1219 => N_1219_5, N_1220 => 
        N_1220_5, BIBUF_COREI2C_0_2_SCL_IO_Y => 
        BIBUF_COREI2C_0_2_SCL_IO_Y, BIBUF_COREI2C_0_2_SDA_IO_Y
         => BIBUF_COREI2C_0_2_SDA_IO_Y, N_1214 => N_1214_3, 
        N_1215 => N_1215_3, N_1216 => N_1216_2, un3_penable_1 => 
        un3_penable_1_0, un105_ens1_1 => un105_ens1_1, N_40 => 
        N_40, un5_penable_1 => un5_penable_1);
    
    BIBUF_COREI2C_0_4_SDA_IO : BIBUF
      port map(PAD => COREI2C_0_4_SDA_IO, D => GND_net_1, E => 
        \COREI2C_0_4_SDAO_i[0]\, Y => BIBUF_COREI2C_0_4_SDA_IO_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity M2sExt_IO_0_IO is

    port( IO_0_Y : out   std_logic_vector(0 to 0);
          PAD_IN : in    std_logic_vector(0 to 0)
        );

end M2sExt_IO_0_IO;

architecture DEF_ARCH of M2sExt_IO_0_IO is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : INBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => PAD_IN(0), Y => IO_0_Y(0));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity M2sExt is

    port( GPIO_IN            : in    std_logic_vector(19 downto 4);
          PAD_IN             : in    std_logic_vector(0 to 0);
          GPIO_OUT           : out   std_logic_vector(2 downto 1);
          USB_ULPI_DATA      : inout std_logic_vector(7 downto 0) := (others => 'Z');
          DEVRST_N           : in    std_logic;
          USB_ULPI_DIR       : in    std_logic;
          USB_ULPI_NXT       : in    std_logic;
          USB_ULPI_XCLK      : in    std_logic;
          USB_RST            : out   std_logic;
          USB_ULPI_STP       : out   std_logic;
          COREI2C_0_0_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_0_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_1_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_1_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_2_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_2_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_3_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_3_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_4_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_4_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_5_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_5_SDA_IO : inout std_logic := 'Z';
          COREI2C_0_6_SCL_IO : inout std_logic := 'Z';
          COREI2C_0_6_SDA_IO : inout std_logic := 'Z'
        );

end M2sExt;

architecture DEF_ARCH of M2sExt is 

  component M2sExt_sb
    port( IO_0_Y             : in    std_logic_vector(0 to 0) := (others => 'U');
          GPIO_IN_c          : in    std_logic_vector(19 downto 4) := (others => 'U');
          GPIO_OUT_c         : out   std_logic_vector(2 downto 1);
          USB_ULPI_DATA      : inout   std_logic_vector(7 downto 0);
          COREI2C_0_6_SDA_IO : inout   std_logic;
          COREI2C_0_6_SCL_IO : inout   std_logic;
          COREI2C_0_5_SDA_IO : inout   std_logic;
          COREI2C_0_5_SCL_IO : inout   std_logic;
          COREI2C_0_4_SDA_IO : inout   std_logic;
          COREI2C_0_4_SCL_IO : inout   std_logic;
          COREI2C_0_3_SDA_IO : inout   std_logic;
          COREI2C_0_3_SCL_IO : inout   std_logic;
          COREI2C_0_2_SDA_IO : inout   std_logic;
          COREI2C_0_2_SCL_IO : inout   std_logic;
          COREI2C_0_1_SDA_IO : inout   std_logic;
          COREI2C_0_1_SCL_IO : inout   std_logic;
          COREI2C_0_0_SDA_IO : inout   std_logic;
          COREI2C_0_0_SCL_IO : inout   std_logic;
          DEVRST_N           : in    std_logic := 'U';
          USB_RST_c          : out   std_logic;
          USB_ULPI_XCLK      : in    std_logic := 'U';
          USB_ULPI_STP       : out   std_logic;
          USB_ULPI_NXT       : in    std_logic := 'U';
          USB_ULPI_DIR       : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component M2sExt_IO_0_IO
    port( IO_0_Y : out   std_logic_vector(0 to 0);
          PAD_IN : in    std_logic_vector(0 to 0) := (others => 'U')
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \IO_0_Y[0]\, VCC_net_1, GND_net_1, \GPIO_IN_c[4]\, 
        \GPIO_IN_c[5]\, \GPIO_IN_c[6]\, \GPIO_IN_c[7]\, 
        \GPIO_IN_c[8]\, \GPIO_IN_c[9]\, \GPIO_IN_c[10]\, 
        \GPIO_IN_c[11]\, \GPIO_IN_c[12]\, \GPIO_IN_c[13]\, 
        \GPIO_IN_c[14]\, \GPIO_IN_c[15]\, \GPIO_IN_c[16]\, 
        \GPIO_IN_c[17]\, \GPIO_IN_c[18]\, \GPIO_IN_c[19]\, 
        \GPIO_OUT_c[1]\, \GPIO_OUT_c[2]\, USB_RST_c : std_logic;

    for all : M2sExt_sb
	Use entity work.M2sExt_sb(DEF_ARCH);
    for all : M2sExt_IO_0_IO
	Use entity work.M2sExt_IO_0_IO(DEF_ARCH);
begin 


    M2sExt_sb_0 : M2sExt_sb
      port map(IO_0_Y(0) => \IO_0_Y[0]\, GPIO_IN_c(19) => 
        \GPIO_IN_c[19]\, GPIO_IN_c(18) => \GPIO_IN_c[18]\, 
        GPIO_IN_c(17) => \GPIO_IN_c[17]\, GPIO_IN_c(16) => 
        \GPIO_IN_c[16]\, GPIO_IN_c(15) => \GPIO_IN_c[15]\, 
        GPIO_IN_c(14) => \GPIO_IN_c[14]\, GPIO_IN_c(13) => 
        \GPIO_IN_c[13]\, GPIO_IN_c(12) => \GPIO_IN_c[12]\, 
        GPIO_IN_c(11) => \GPIO_IN_c[11]\, GPIO_IN_c(10) => 
        \GPIO_IN_c[10]\, GPIO_IN_c(9) => \GPIO_IN_c[9]\, 
        GPIO_IN_c(8) => \GPIO_IN_c[8]\, GPIO_IN_c(7) => 
        \GPIO_IN_c[7]\, GPIO_IN_c(6) => \GPIO_IN_c[6]\, 
        GPIO_IN_c(5) => \GPIO_IN_c[5]\, GPIO_IN_c(4) => 
        \GPIO_IN_c[4]\, GPIO_OUT_c(2) => \GPIO_OUT_c[2]\, 
        GPIO_OUT_c(1) => \GPIO_OUT_c[1]\, USB_ULPI_DATA(7) => 
        USB_ULPI_DATA(7), USB_ULPI_DATA(6) => USB_ULPI_DATA(6), 
        USB_ULPI_DATA(5) => USB_ULPI_DATA(5), USB_ULPI_DATA(4)
         => USB_ULPI_DATA(4), USB_ULPI_DATA(3) => 
        USB_ULPI_DATA(3), USB_ULPI_DATA(2) => USB_ULPI_DATA(2), 
        USB_ULPI_DATA(1) => USB_ULPI_DATA(1), USB_ULPI_DATA(0)
         => USB_ULPI_DATA(0), COREI2C_0_6_SDA_IO => 
        COREI2C_0_6_SDA_IO, COREI2C_0_6_SCL_IO => 
        COREI2C_0_6_SCL_IO, COREI2C_0_5_SDA_IO => 
        COREI2C_0_5_SDA_IO, COREI2C_0_5_SCL_IO => 
        COREI2C_0_5_SCL_IO, COREI2C_0_4_SDA_IO => 
        COREI2C_0_4_SDA_IO, COREI2C_0_4_SCL_IO => 
        COREI2C_0_4_SCL_IO, COREI2C_0_3_SDA_IO => 
        COREI2C_0_3_SDA_IO, COREI2C_0_3_SCL_IO => 
        COREI2C_0_3_SCL_IO, COREI2C_0_2_SDA_IO => 
        COREI2C_0_2_SDA_IO, COREI2C_0_2_SCL_IO => 
        COREI2C_0_2_SCL_IO, COREI2C_0_1_SDA_IO => 
        COREI2C_0_1_SDA_IO, COREI2C_0_1_SCL_IO => 
        COREI2C_0_1_SCL_IO, COREI2C_0_0_SDA_IO => 
        COREI2C_0_0_SDA_IO, COREI2C_0_0_SCL_IO => 
        COREI2C_0_0_SCL_IO, DEVRST_N => DEVRST_N, USB_RST_c => 
        USB_RST_c, USB_ULPI_XCLK => USB_ULPI_XCLK, USB_ULPI_STP
         => USB_ULPI_STP, USB_ULPI_NXT => USB_ULPI_NXT, 
        USB_ULPI_DIR => USB_ULPI_DIR);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \GPIO_IN_ibuf[15]\ : INBUF
      port map(PAD => GPIO_IN(15), Y => \GPIO_IN_c[15]\);
    
    \GPIO_IN_ibuf[12]\ : INBUF
      port map(PAD => GPIO_IN(12), Y => \GPIO_IN_c[12]\);
    
    IO_0 : M2sExt_IO_0_IO
      port map(IO_0_Y(0) => \IO_0_Y[0]\, PAD_IN(0) => PAD_IN(0));
    
    \GPIO_IN_ibuf[6]\ : INBUF
      port map(PAD => GPIO_IN(6), Y => \GPIO_IN_c[6]\);
    
    \GPIO_IN_ibuf[16]\ : INBUF
      port map(PAD => GPIO_IN(16), Y => \GPIO_IN_c[16]\);
    
    \GPIO_OUT_obuf[2]\ : OUTBUF
      port map(D => \GPIO_OUT_c[2]\, PAD => GPIO_OUT(2));
    
    \GPIO_OUT_obuf[1]\ : OUTBUF
      port map(D => \GPIO_OUT_c[1]\, PAD => GPIO_OUT(1));
    
    \GPIO_IN_ibuf[4]\ : INBUF
      port map(PAD => GPIO_IN(4), Y => \GPIO_IN_c[4]\);
    
    \GPIO_IN_ibuf[8]\ : INBUF
      port map(PAD => GPIO_IN(8), Y => \GPIO_IN_c[8]\);
    
    \GPIO_IN_ibuf[19]\ : INBUF
      port map(PAD => GPIO_IN(19), Y => \GPIO_IN_c[19]\);
    
    \GPIO_IN_ibuf[17]\ : INBUF
      port map(PAD => GPIO_IN(17), Y => \GPIO_IN_c[17]\);
    
    \GPIO_IN_ibuf[14]\ : INBUF
      port map(PAD => GPIO_IN(14), Y => \GPIO_IN_c[14]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GPIO_IN_ibuf[7]\ : INBUF
      port map(PAD => GPIO_IN(7), Y => \GPIO_IN_c[7]\);
    
    \GPIO_IN_ibuf[5]\ : INBUF
      port map(PAD => GPIO_IN(5), Y => \GPIO_IN_c[5]\);
    
    \GPIO_IN_ibuf[18]\ : INBUF
      port map(PAD => GPIO_IN(18), Y => \GPIO_IN_c[18]\);
    
    \GPIO_IN_ibuf[9]\ : INBUF
      port map(PAD => GPIO_IN(9), Y => \GPIO_IN_c[9]\);
    
    \GPIO_IN_ibuf[11]\ : INBUF
      port map(PAD => GPIO_IN(11), Y => \GPIO_IN_c[11]\);
    
    \GPIO_IN_ibuf[10]\ : INBUF
      port map(PAD => GPIO_IN(10), Y => \GPIO_IN_c[10]\);
    
    USB_RST_obuf : OUTBUF
      port map(D => USB_RST_c, PAD => USB_RST);
    
    \GPIO_IN_ibuf[13]\ : INBUF
      port map(PAD => GPIO_IN(13), Y => \GPIO_IN_c[13]\);
    

end DEF_ARCH; 
